        nop(32);
        activate(2, 329);
        nop(6);
        activate(1, 1587);
        nop(5);
        read(2, 95, 0, 0);
        nop(1);
        activate(6, 394);
        nop(3);
        read(2, 95, 0, 0);
        nop(3);
        activate(7, 447);
        nop(1);
        read(1, 5, 0, 0);
        nop(4);
        read(1, 5, 0, 0);
        nop(4);
        read(1, 5, 0, 0);
        nop(4);
        read(1, 5, 0, 0);
        nop(4);
        read(2, 95, 0, 0);
        nop(4);
        read(7, 73, 0, 0);
        nop(4);
        read(7, 73, 0, 0);
        nop(4);
        read(7, 73, 0, 0);
        nop(4);
        read(7, 73, 0, 0);
        nop(4);
        read(7, 73, 0, 0);
        nop(4);
        read(1, 6, 0, 0);
        nop(4);
        read(1, 6, 0, 0);
        nop(4);
        read(2, 95, 0, 0);
        nop(4);
        read(7, 73, 0, 0);
        nop(4);
        read(7, 73, 0, 0);
        nop(4);
        read(7, 73, 0, 0);
        nop(4);
        read(1, 6, 0, 0);
        nop(4);
        read(1, 6, 0, 0);
        nop(2);
        activate(0, 494);
        nop(2);
        read(1, 6, 0, 0);
        nop(4);
        read(2, 95, 0, 0);
        nop(4);
        read(1, 6, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(2);
        read(0, 58, 0, 0);
        nop(4);
        read(0, 58, 0, 0);
        nop(4);
        read(0, 58, 0, 0);
        nop(2);
        activate(2, 329);
        nop(2);
        read(1, 6, 0, 0);
        nop(4);
        read(0, 58, 0, 0);
        nop(4);
        read(0, 58, 0, 0);
        nop(4);
        read(0, 58, 0, 0);
        nop(4);
        read(0, 58, 0, 0);
        nop(4);
        read(0, 58, 0, 0);
        nop(4);
        read(1, 6, 0, 0);
        nop(4);
        read(1, 7, 0, 0);
        nop(4);
        read(1, 7, 0, 0);
        nop(4);
        read(2, 96, 0, 0);
        nop(4);
        read(1, 7, 0, 0);
        nop(4);
        read(1, 7, 0, 0);
        nop(4);
        read(2, 96, 0, 0);
        nop(4);
        read(2, 96, 0, 0);
        nop(4);
        read(2, 96, 0, 0);
        nop(4);
        read(1, 7, 0, 0);
        nop(4);
        read(1, 7, 0, 0);
        nop(4);
        read(2, 96, 0, 0);
        nop(4);
        read(1, 7, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(2);
        read(1, 7, 0, 0);
        nop(4);
        read(1, 8, 0, 0);
        nop(4);
        read(1, 8, 0, 0);
        nop(2);
        activate(2, 329);
        nop(2);
        read(1, 8, 0, 0);
        nop(4);
        read(1, 8, 0, 0);
        nop(4);
        read(1, 8, 0, 0);
        nop(4);
        read(1, 8, 0, 0);
        nop(2);
        precharge(7, 0);
        nop(2);
        read(1, 8, 0, 0);
        nop(4);
        read(1, 8, 0, 0);
        nop(4);
        read(2, 95, 0, 0);
        nop(2);
        activate(7, 447);
        nop(2);
        read(2, 95, 0, 0);
        nop(2);
        precharge(0, 0);
        nop(2);
        read(2, 95, 0, 0);
        nop(4);
        read(2, 94, 0, 0);
        nop(4);
        read(7, 80, 0, 0);
        nop(2);
        activate(0, 321);
        nop(2);
        read(2, 94, 0, 0);
        nop(4);
        read(7, 80, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(2);
        read(7, 80, 0, 0);
        nop(4);
        read(7, 80, 0, 0);
        nop(4);
        read(0, 42, 0, 0);
        nop(2);
        activate(2, 329);
        nop(2);
        read(0, 42, 0, 0);
        nop(4);
        read(0, 42, 0, 0);
        nop(1);
        activate(3, 2026);
        nop(3);
        read(0, 42, 0, 0);
        nop(4);
        read(0, 42, 0, 0);
        nop(4);
        read(0, 42, 0, 0);
        nop(4);
        read(0, 42, 0, 0);
        nop(4);
        read(0, 42, 0, 0);
        nop(4);
        read(2, 96, 0, 0);
        nop(4);
        read(2, 96, 0, 0);
        nop(4);
        read(2, 96, 0, 0);
        nop(4);
        read(3, 108, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(7);
        write(6, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(6, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(1);
        activate(2, 329);
        nop(3);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(17);
        read(2, 94, 0, 0);
        nop(2);
        precharge(6, 0);
        nop(2);
        read(2, 94, 0, 0);
        nop(4);
        read(3, 108, 0, 0);
        nop(4);
        read(2, 94, 0, 0);
        nop(2);
        activate(6, 421);
        nop(2);
        read(2, 94, 0, 0);
        nop(4);
        read(2, 94, 0, 0);
        nop(4);
        read(2, 94, 0, 0);
        nop(4);
        read(6, 109, 0, 0);
        nop(4);
        read(6, 109, 0, 0);
        nop(4);
        read(6, 109, 0, 0);
        nop(4);
        read(6, 109, 0, 0);
        nop(4);
        read(6, 109, 0, 0);
        nop(6);
        precharge(6, 0);
        nop(3);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(9);
        activate(6, 406);
        nop(8);
        read(3, 108, 0, 0);
        nop(4);
        read(6, 62, 0, 0);
        nop(4);
        read(6, 62, 0, 0);
        nop(4);
        read(6, 62, 0, 0);
        nop(4);
        read(6, 62, 0, 0);
        nop(4);
        read(6, 62, 0, 0);
        nop(6);
        precharge(6, 0);
        nop(3);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(9);
        activate(6, 421);
        nop(8);
        read(3, 108, 0, 0);
        nop(4);
        read(6, 109, 0, 0);
        nop(4);
        read(6, 109, 0, 0);
        nop(4);
        read(6, 109, 0, 0);
        nop(4);
        read(0, 43, 0, 0);
        nop(4);
        read(0, 43, 0, 0);
        nop(1);
        precharge(6, 0);
        nop(3);
        read(0, 43, 0, 0);
        nop(4);
        read(0, 43, 0, 0);
        nop(4);
        read(0, 43, 0, 0);
        nop(1);
        activate(6, 406);
        nop(3);
        read(0, 43, 0, 0);
        nop(4);
        read(0, 43, 0, 0);
        nop(4);
        read(0, 43, 0, 0);
        nop(4);
        read(6, 62, 0, 0);
        nop(4);
        read(6, 62, 0, 0);
        nop(4);
        read(6, 62, 0, 0);
        nop(9);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(505);
        read(0, 44, 0, 0);
        nop(4);
        read(0, 44, 0, 0);
        nop(1);
        activate(4, 393);
        nop(3);
        read(0, 44, 0, 0);
        nop(4);
        read(0, 44, 0, 0);
        nop(4);
        read(4, 70, 0, 0);
        nop(4);
        read(4, 70, 0, 0);
        nop(4);
        read(4, 70, 0, 0);
        nop(4);
        read(4, 70, 0, 0);
        nop(4);
        read(0, 44, 0, 0);
        nop(4);
        read(0, 44, 0, 0);
        nop(4);
        read(0, 44, 0, 0);
        nop(4);
        read(0, 44, 0, 0);
        nop(4);
        read(3, 108, 0, 0);
        nop(9);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(115);
        read(3, 108, 0, 0);
        nop(9);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(17);
        read(3, 108, 0, 0);
        nop(9);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(120);
        read(3, 108, 0, 0);
        nop(6);
        precharge(2, 0);
        nop(3);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(9);
        activate(2, 423);
        nop(10);
        precharge(7, 0);
        nop(1);
        read(2, 54, 0, 0);
        nop(2);
        precharge(4, 0);
        nop(2);
        read(2, 54, 0, 0);
        nop(3);
        precharge(0, 0);
        nop(1);
        read(2, 54, 0, 0);
        nop(3);
        activate(7, 1560);
        nop(1);
        read(2, 54, 0, 0);
        nop(4);
        read(2, 54, 0, 0);
        nop(1);
        activate(4, 1887);
        nop(5);
        read(7, 64, 0, 0);
        nop(1);
        activate(0, 265);
        nop(1);
        precharge(2, 0);
        nop(2);
        read(7, 64, 0, 0);
        nop(4);
        read(4, 4, 0, 0);
        nop(4);
        read(4, 4, 0, 0);
        nop(2);
        activate(2, 481);
        nop(2);
        read(4, 4, 0, 0);
        nop(4);
        read(7, 64, 0, 0);
        nop(4);
        read(7, 64, 0, 0);
        nop(4);
        read(0, 20, 0, 0);
        nop(4);
        read(0, 20, 0, 0);
        nop(4);
        read(4, 4, 0, 0);
        nop(4);
        read(4, 4, 0, 0);
        nop(4);
        read(0, 20, 0, 0);
        nop(2);
        precharge(4, 0);
        nop(2);
        read(0, 20, 0, 0);
        nop(4);
        read(0, 20, 0, 0);
        nop(6);
        precharge(0, 0);
        nop(1);
        activate(4, 447);
        nop(2);
        write(2, 54, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(2, 54, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(2, 54, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(1);
        activate(0, 321);
        nop(3);
        write(2, 54, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(17);
        read(0, 45, 0, 0);
        nop(4);
        read(0, 45, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(2);
        read(4, 95, 0, 0);
        nop(4);
        read(4, 95, 0, 0);
        nop(4);
        read(4, 95, 0, 0);
        nop(2);
        activate(2, 423);
        nop(2);
        read(0, 45, 0, 0);
        nop(4);
        read(0, 45, 0, 0);
        nop(4);
        read(0, 45, 0, 0);
        nop(4);
        read(2, 54, 0, 0);
        nop(2);
        precharge(0, 0);
        nop(2);
        read(2, 54, 0, 0);
        nop(4);
        read(4, 95, 0, 0);
        nop(4);
        read(2, 54, 0, 0);
        nop(2);
        activate(0, 265);
        nop(1);
        precharge(4, 0);
        nop(1);
        read(2, 55, 0, 0);
        nop(4);
        read(2, 55, 0, 0);
        nop(5);
        read(0, 20, 0, 0);
        nop(1);
        precharge(2, 0);
        nop(1);
        activate(4, 1887);
        nop(2);
        read(0, 20, 0, 0);
        nop(4);
        read(0, 20, 0, 0);
        nop(5);
        activate(2, 329);
        nop(1);
        read(4, 4, 0, 0);
        nop(3);
        precharge(0, 0);
        nop(1);
        read(4, 4, 0, 0);
        nop(4);
        read(4, 4, 0, 0);
        nop(4);
        read(2, 122, 0, 0);
        nop(3);
        activate(0, 321);
        nop(1);
        read(2, 122, 0, 0);
        nop(4);
        read(2, 122, 0, 0);
        nop(4);
        read(2, 122, 0, 0);
        nop(2);
        precharge(4, 0);
        nop(2);
        read(2, 122, 0, 0);
        nop(4);
        read(0, 45, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(2);
        read(0, 45, 0, 0);
        nop(2);
        activate(5, 450);
        nop(2);
        read(0, 45, 0, 0);
        nop(4);
        activate(4, 508);
        nop(5);
        read(5, 74, 0, 0);
        nop(1);
        activate(2, 423);
        nop(3);
        read(5, 74, 0, 0);
        nop(4);
        read(4, 19, 0, 0);
        nop(4);
        read(4, 19, 0, 0);
        nop(4);
        read(5, 74, 0, 0);
        nop(4);
        read(2, 55, 0, 0);
        nop(4);
        read(2, 55, 0, 0);
        nop(4);
        read(2, 55, 0, 0);
        nop(4);
        read(2, 55, 0, 0);
        nop(4);
        read(2, 55, 0, 0);
        nop(4);
        read(4, 19, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(2);
        read(5, 74, 0, 0);
        nop(4);
        read(4, 19, 0, 0);
        nop(4);
        read(5, 74, 0, 0);
        nop(2);
        activate(2, 329);
        nop(4);
        precharge(5, 0);
        nop(7);
        read(2, 122, 0, 0);
        nop(4);
        read(2, 122, 0, 0);
        nop(1);
        activate(5, 503);
        nop(3);
        read(2, 122, 0, 0);
        nop(4);
        read(2, 123, 0, 0);
        nop(4);
        read(2, 123, 0, 0);
        nop(6);
        precharge(2, 0);
        nop(3);
        write(5, 74, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(5, 74, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(5, 74, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(1);
        activate(2, 423);
        nop(3);
        write(5, 74, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(17);
        read(2, 55, 0, 0);
        nop(6);
        precharge(5, 0);
        nop(2);
        precharge(2, 0);
        nop(10);
        activate(5, 450);
        nop(6);
        activate(2, 329);
        nop(5);
        read(5, 74, 0, 0);
        nop(4);
        read(5, 74, 0, 0);
        nop(4);
        read(5, 74, 0, 0);
        nop(4);
        read(2, 123, 0, 0);
        nop(4);
        read(2, 123, 0, 0);
        nop(1);
        precharge(5, 0);
        nop(3);
        read(2, 124, 0, 0);
        nop(4);
        read(2, 124, 0, 0);
        nop(4);
        read(2, 124, 0, 0);
        nop(1);
        activate(5, 441);
        nop(5);
        precharge(2, 0);
        nop(6);
        read(5, 84, 0, 0);
        nop(4);
        read(5, 84, 0, 0);
        nop(2);
        activate(2, 399);
        nop(2);
        read(5, 84, 0, 0);
        nop(4);
        read(5, 84, 0, 0);
        nop(6);
        precharge(5, 0);
        nop(3);
        write(2, 125, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(2, 125, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(2, 125, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(1);
        activate(5, 452);
        nop(3);
        write(2, 125, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(2);
        precharge(4, 0);
        nop(12);
        activate(4, 476);
        nop(3);
        read(5, 84, 0, 0);
        nop(4);
        read(5, 84, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(2);
        read(4, 88, 0, 0);
        nop(4);
        read(4, 88, 0, 0);
        nop(4);
        read(4, 88, 0, 0);
        nop(2);
        activate(2, 329);
        nop(2);
        read(4, 88, 0, 0);
        nop(4);
        read(4, 88, 0, 0);
        nop(4);
        read(4, 88, 0, 0);
        nop(4);
        read(5, 84, 0, 0);
        nop(2);
        precharge(4, 0);
        nop(2);
        read(2, 124, 0, 0);
        nop(4);
        read(2, 125, 0, 0);
        nop(4);
        read(2, 125, 0, 0);
        nop(2);
        activate(4, 508);
        nop(2);
        read(5, 84, 0, 0);
        nop(4);
        read(2, 125, 0, 0);
        nop(2);
        precharge(5, 0);
        nop(2);
        read(2, 125, 0, 0);
        nop(2);
        precharge(6, 0);
        nop(2);
        read(2, 125, 0, 0);
        nop(4);
        read(2, 125, 0, 0);
        nop(2);
        activate(5, 363);
        nop(2);
        read(4, 20, 0, 0);
        nop(2);
        precharge(7, 0);
        nop(2);
        activate(6, 492);
        nop(1);
        read(2, 125, 0, 0);
        nop(4);
        read(2, 125, 0, 0);
        nop(4);
        read(4, 20, 0, 0);
        nop(1);
        activate(7, 501);
        nop(3);
        read(4, 20, 0, 0);
        nop(2);
        precharge(0, 0);
        nop(2);
        read(4, 20, 0, 0);
        nop(4);
        read(6, 17, 0, 0);
        nop(4);
        read(6, 17, 0, 0);
        nop(2);
        activate(0, 406);
        nop(1);
        precharge(3, 0);
        nop(1);
        read(4, 20, 0, 0);
        nop(4);
        read(6, 17, 0, 0);
        nop(2);
        precharge(4, 0);
        nop(2);
        read(6, 17, 0, 0);
        nop(3);
        activate(3, 510);
        nop(1);
        read(7, 94, 0, 0);
        nop(4);
        read(7, 94, 0, 0);
        nop(2);
        activate(4, 476);
        nop(2);
        read(7, 94, 0, 0);
        nop(4);
        read(3, 5, 0, 0);
        nop(4);
        read(3, 5, 0, 0);
        nop(4);
        read(4, 88, 0, 0);
        nop(4);
        read(7, 94, 0, 0);
        nop(4);
        read(0, 38, 0, 0);
        nop(4);
        read(0, 38, 0, 0);
        nop(4);
        read(0, 38, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(2);
        read(3, 5, 0, 0);
        nop(4);
        read(3, 5, 0, 0);
        nop(4);
        read(4, 88, 0, 0);
        nop(2);
        activate(2, 503);
        nop(2);
        read(0, 38, 0, 0);
        nop(2);
        precharge(4, 0);
        nop(2);
        read(3, 5, 0, 0);
        nop(5);
        read(2, 65, 0, 0);
        nop(1);
        precharge(3, 0);
        nop(3);
        read(2, 65, 0, 0);
        nop(1);
        activate(4, 508);
        nop(3);
        read(2, 65, 0, 0);
        nop(4);
        read(2, 65, 0, 0);
        nop(1);
        activate(3, 510);
        nop(3);
        read(4, 20, 0, 0);
        nop(4);
        read(4, 20, 0, 0);
        nop(4);
        read(3, 85, 0, 0);
        nop(4);
        read(3, 85, 0, 0);
        nop(4);
        read(4, 20, 0, 0);
        nop(4);
        read(3, 85, 0, 0);
        nop(4);
        read(3, 85, 0, 0);
        nop(6);
        precharge(3, 0);
        nop(3);
        write(5, 84, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(5, 84, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(5, 84, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(1);
        activate(3, 510);
        nop(3);
        write(5, 84, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(17);
        read(3, 5, 0, 0);
        nop(4);
        read(3, 5, 0, 0);
        nop(2);
        precharge(5, 0);
        nop(2);
        read(3, 5, 0, 0);
        nop(4);
        read(4, 21, 0, 0);
        nop(2);
        precharge(3, 0);
        nop(2);
        read(4, 21, 0, 0);
        nop(2);
        activate(5, 452);
        nop(2);
        read(4, 21, 0, 0);
        nop(4);
        read(4, 21, 0, 0);
        nop(2);
        activate(3, 440);
        nop(2);
        read(4, 21, 0, 0);
        nop(4);
        read(4, 21, 0, 0);
        nop(2);
        precharge(7, 0);
        nop(2);
        read(4, 21, 0, 0);
        nop(4);
        read(4, 21, 0, 0);
        nop(4);
        read(5, 66, 0, 0);
        nop(2);
        activate(7, 516);
        nop(2);
        read(3, 11, 0, 0);
        nop(4);
        read(3, 11, 0, 0);
        nop(4);
        read(3, 11, 0, 0);
        nop(4);
        read(3, 11, 0, 0);
        nop(4);
        read(3, 11, 0, 0);
        nop(2);
        precharge(4, 0);
        nop(2);
        read(5, 66, 0, 0);
        nop(2);
        precharge(3, 0);
        nop(2);
        read(7, 13, 0, 0);
        nop(4);
        read(5, 66, 0, 0);
        nop(2);
        activate(4, 393);
        nop(2);
        read(5, 66, 0, 0);
        nop(4);
        activate(3, 440);
        nop(1);
        read(7, 13, 0, 0);
        nop(1);
        precharge(5, 0);
        nop(3);
        read(7, 13, 0, 0);
        nop(4);
        read(7, 13, 0, 0);
        nop(2);
        precharge(0, 0);
        nop(2);
        read(3, 29, 0, 0);
        nop(1);
        activate(5, 933);
        nop(3);
        read(3, 29, 0, 0);
        nop(4);
        read(4, 75, 0, 0);
        nop(2);
        activate(0, 321);
        nop(2);
        read(7, 13, 0, 0);
        nop(4);
        read(7, 13, 0, 0);
        nop(4);
        read(3, 29, 0, 0);
        nop(4);
        read(3, 29, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(2);
        read(3, 29, 0, 0);
        nop(4);
        read(4, 75, 0, 0);
        nop(2);
        precharge(3, 0);
        nop(2);
        read(7, 13, 0, 0);
        nop(2);
        activate(2, 329);
        nop(2);
        read(0, 46, 0, 0);
        nop(4);
        read(4, 75, 0, 0);
        nop(2);
        activate(3, 440);
        nop(2);
        read(4, 75, 0, 0);
        nop(4);
        read(4, 75, 0, 0);
        nop(4);
        read(7, 13, 0, 0);
        nop(4);
        read(0, 46, 0, 0);
        nop(4);
        read(0, 46, 0, 0);
        nop(4);
        read(0, 46, 0, 0);
        nop(4);
        read(2, 127, 0, 0);
        nop(4);
        read(2, 127, 0, 0);
        nop(4);
        read(3, 11, 0, 0);
        nop(4);
        read(4, 75, 0, 0);
        nop(4);
        read(0, 46, 0, 0);
        nop(4);
        read(0, 46, 0, 0);
        nop(4);
        read(0, 46, 0, 0);
        nop(4);
        read(0, 46, 0, 0);
        nop(4);
        read(2, 127, 0, 0);
        nop(4);
        read(2, 127, 0, 0);
        nop(4);
        read(3, 11, 0, 0);
        nop(4);
        read(4, 75, 0, 0);
        nop(4);
        read(2, 127, 0, 0);
        nop(4);
        read(2, 127, 0, 0);
        nop(4);
        read(2, 127, 0, 0);
        nop(4);
        read(2, 127, 0, 0);
        nop(4);
        read(3, 11, 0, 0);
        nop(4);
        read(4, 75, 0, 0);
        nop(2);
        precharge(3, 0);
        nop(7);
        write(5, 66, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(5, 66, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(1);
        activate(3, 440);
        nop(3);
        write(5, 66, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(5, 66, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(17);
        read(3, 29, 0, 0);
        nop(4);
        read(3, 29, 0, 0);
        nop(2);
        precharge(5, 0);
        nop(2);
        read(3, 29, 0, 0);
        nop(10);
        activate(5, 1831);
        nop(11);
        read(5, 22, 0, 0);
        nop(4);
        read(5, 22, 0, 0);
        nop(4);
        read(5, 22, 0, 0);
        nop(4);
        read(5, 22, 0, 0);
        nop(4);
        read(5, 22, 0, 0);
        nop(6);
        precharge(5, 0);
        nop(12);
        activate(5, 329);
        nop(11);
        read(5, 65, 0, 0);
        nop(4);
        read(5, 65, 0, 0);
        nop(4);
        read(5, 65, 0, 0);
        nop(4);
        read(5, 65, 0, 0);
        nop(4);
        read(5, 65, 0, 0);
        nop(6);
        precharge(5, 0);
        nop(12);
        activate(5, 1831);
        nop(11);
        read(5, 22, 0, 0);
        nop(4);
        read(5, 22, 0, 0);
        nop(4);
        read(5, 22, 0, 0);
        nop(9);
        precharge(5, 0);
        nop(12);
        activate(5, 329);
        nop(11);
        read(5, 65, 0, 0);
        nop(4);
        read(5, 65, 0, 0);
        nop(4);
        read(5, 65, 0, 0);
        nop(4);
        read(5, 66, 0, 0);
        nop(4);
        read(5, 66, 0, 0);
        nop(4);
        read(5, 66, 0, 0);
        nop(4);
        read(5, 66, 0, 0);
        nop(4);
        read(5, 66, 0, 0);
        nop(4);
        read(5, 66, 0, 0);
        nop(4);
        read(5, 66, 0, 0);
        nop(4);
        read(5, 66, 0, 0);
        nop(4);
        read(5, 67, 0, 0);
        nop(4);
        read(5, 67, 0, 0);
        nop(4);
        read(5, 67, 0, 0);
        nop(4);
        read(5, 67, 0, 0);
        nop(4);
        read(5, 67, 0, 0);
        nop(4);
        read(5, 67, 0, 0);
        nop(4);
        read(5, 67, 0, 0);
        nop(4);
        read(5, 67, 0, 0);
        nop(2);
        precharge(7, 0);
        nop(2);
        read(5, 68, 0, 0);
        nop(4);
        read(5, 68, 0, 0);
        nop(4);
        read(5, 68, 0, 0);
        nop(2);
        precharge(3, 0);
        nop(1);
        activate(7, 513);
        nop(1);
        read(5, 68, 0, 0);
        nop(4);
        read(5, 68, 0, 0);
        nop(4);
        read(5, 68, 0, 0);
        nop(2);
        activate(3, 2026);
        nop(2);
        read(7, 72, 0, 0);
        nop(4);
        read(7, 72, 0, 0);
        nop(4);
        read(5, 68, 0, 0);
        nop(4);
        read(3, 108, 0, 0);
        nop(4);
        read(5, 68, 0, 0);
        nop(4);
        read(7, 72, 0, 0);
        nop(2);
        precharge(5, 0);
        nop(2);
        read(7, 72, 0, 0);
        nop(9);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(1);
        activate(5, 422);
        nop(16);
        read(3, 108, 0, 0);
        nop(4);
        read(5, 70, 0, 0);
        nop(4);
        read(5, 70, 0, 0);
        nop(4);
        read(5, 70, 0, 0);
        nop(4);
        read(5, 70, 0, 0);
        nop(2);
        precharge(0, 0);
        nop(2);
        read(5, 70, 0, 0);
        nop(6);
        precharge(5, 0);
        nop(3);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(1);
        activate(0, 321);
        nop(8);
        activate(5, 329);
        nop(8);
        read(3, 108, 0, 0);
        nop(4);
        read(5, 70, 0, 0);
        nop(4);
        read(5, 70, 0, 0);
        nop(4);
        read(0, 48, 0, 0);
        nop(4);
        read(0, 48, 0, 0);
        nop(4);
        read(0, 48, 0, 0);
        nop(4);
        read(5, 70, 0, 0);
        nop(4);
        read(5, 70, 0, 0);
        nop(4);
        read(5, 70, 0, 0);
        nop(4);
        read(0, 48, 0, 0);
        nop(2);
        precharge(5, 0);
        nop(2);
        read(0, 49, 0, 0);
        nop(4);
        read(0, 49, 0, 0);
        nop(4);
        read(0, 49, 0, 0);
        nop(2);
        activate(5, 422);
        nop(2);
        read(0, 49, 0, 0);
        nop(4);
        read(0, 49, 0, 0);
        nop(4);
        read(0, 49, 0, 0);
        nop(4);
        read(5, 70, 0, 0);
        nop(4);
        read(0, 49, 0, 0);
        nop(4);
        read(0, 49, 0, 0);
        nop(4);
        read(0, 50, 0, 0);
        nop(4);
        read(5, 70, 0, 0);
        nop(4);
        read(5, 70, 0, 0);
        nop(4);
        read(0, 50, 0, 0);
        nop(2);
        precharge(5, 0);
        nop(2);
        read(0, 50, 0, 0);
        nop(4);
        read(0, 50, 0, 0);
        nop(4);
        read(0, 50, 0, 0);
        nop(2);
        activate(5, 329);
        nop(2);
        read(0, 50, 0, 0);
        nop(4);
        read(0, 50, 0, 0);
        nop(4);
        read(0, 50, 0, 0);
        nop(4);
        read(5, 70, 0, 0);
        nop(4);
        read(5, 70, 0, 0);
        nop(4);
        read(5, 70, 0, 0);
        nop(4);
        read(5, 71, 0, 0);
        nop(4);
        read(5, 71, 0, 0);
        nop(6);
        precharge(5, 0);
        nop(3);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(9);
        activate(5, 329);
        nop(8);
        read(3, 108, 0, 0);
        nop(4);
        read(5, 80, 0, 0);
        nop(4);
        read(5, 80, 0, 0);
        nop(4);
        read(5, 80, 0, 0);
        nop(4);
        read(5, 80, 0, 0);
        nop(4);
        read(5, 81, 0, 0);
        nop(6);
        precharge(5, 0);
        nop(3);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(9);
        activate(5, 329);
        nop(11);
        read(5, 71, 0, 0);
        nop(4);
        read(5, 71, 0, 0);
        nop(4);
        read(5, 71, 0, 0);
        nop(4);
        read(5, 71, 0, 0);
        nop(4);
        read(5, 71, 0, 0);
        nop(6);
        precharge(5, 0);
        nop(12);
        activate(5, 329);
        nop(11);
        read(5, 81, 0, 0);
        nop(4);
        read(5, 81, 0, 0);
        nop(4);
        read(5, 81, 0, 0);
        nop(4);
        read(5, 82, 0, 0);
        nop(4);
        read(5, 82, 0, 0);
        nop(6);
        precharge(5, 0);
        nop(12);
        activate(5, 329);
        nop(11);
        read(5, 71, 0, 0);
        nop(4);
        read(5, 72, 0, 0);
        nop(4);
        read(5, 72, 0, 0);
        nop(4);
        read(5, 72, 0, 0);
        nop(4);
        read(5, 72, 0, 0);
        nop(6);
        precharge(5, 0);
        nop(12);
        activate(5, 329);
        nop(11);
        read(5, 82, 0, 0);
        nop(4);
        read(5, 82, 0, 0);
        nop(4);
        read(5, 82, 0, 0);
        nop(4);
        read(5, 82, 0, 0);
        nop(4);
        read(5, 82, 0, 0);
        nop(6);
        precharge(5, 0);
        nop(12);
        activate(5, 329);
        nop(11);
        read(5, 72, 0, 0);
        nop(4);
        read(5, 72, 0, 0);
        nop(4);
        read(5, 72, 0, 0);
        nop(4);
        read(5, 72, 0, 0);
        nop(4);
        read(5, 79, 0, 0);
        nop(2);
        precharge(0, 0);
        nop(4);
        precharge(5, 0);
        nop(8);
        activate(0, 406);
        nop(6);
        activate(5, 329);
        nop(5);
        read(0, 36, 0, 0);
        nop(4);
        read(0, 36, 0, 0);
        nop(4);
        read(5, 82, 0, 0);
        nop(4);
        read(5, 84, 0, 0);
        nop(4);
        read(0, 36, 0, 0);
        nop(4);
        read(0, 36, 0, 0);
        nop(4);
        read(5, 84, 0, 0);
        nop(4);
        read(5, 84, 0, 0);
        nop(4);
        read(5, 84, 0, 0);
        nop(6);
        precharge(5, 0);
        nop(12);
        activate(5, 329);
        nop(11);
        read(5, 79, 0, 0);
        nop(4);
        read(5, 79, 0, 0);
        nop(4);
        read(5, 79, 0, 0);
        nop(4);
        read(5, 79, 0, 0);
        nop(4);
        read(5, 79, 0, 0);
        nop(6);
        precharge(5, 0);
        nop(12);
        activate(5, 509);
        nop(11);
        write(5, 82, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(5, 82, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(5, 82, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(5, 82, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(5, 82, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(17);
        read(3, 108, 0, 0);
        nop(6);
        precharge(5, 0);
        nop(3);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(9);
        activate(5, 329);
        nop(8);
        read(3, 108, 0, 0);
        nop(4);
        read(5, 79, 0, 0);
        nop(2);
        precharge(0, 0);
        nop(2);
        read(5, 79, 0, 0);
        nop(9);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(1);
        activate(0, 321);
        nop(2);
        precharge(5, 0);
        nop(12);
        activate(5, 509);
        nop(2);
        read(0, 52, 0, 0);
        nop(4);
        read(0, 52, 0, 0);
        nop(4);
        read(0, 52, 0, 0);
        nop(4);
        read(0, 52, 0, 0);
        nop(4);
        read(3, 108, 0, 0);
        nop(4);
        read(0, 53, 0, 0);
        nop(4);
        read(0, 53, 0, 0);
        nop(4);
        read(0, 53, 0, 0);
        nop(4);
        read(0, 53, 0, 0);
        nop(4);
        read(0, 53, 0, 0);
        nop(4);
        read(0, 53, 0, 0);
        nop(4);
        read(0, 53, 0, 0);
        nop(4);
        read(0, 53, 0, 0);
        nop(4);
        read(0, 54, 0, 0);
        nop(4);
        read(0, 54, 0, 0);
        nop(4);
        read(0, 54, 0, 0);
        nop(4);
        read(0, 54, 0, 0);
        nop(4);
        read(0, 54, 0, 0);
        nop(4);
        read(0, 54, 0, 0);
        nop(4);
        read(0, 54, 0, 0);
        nop(4);
        read(0, 54, 0, 0);
        nop(9);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(5, 82, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(5, 82, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(5, 82, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(17);
        read(3, 108, 0, 0);
        nop(4);
        read(0, 55, 0, 0);
        nop(2);
        precharge(5, 0);
        nop(2);
        read(0, 55, 0, 0);
        nop(4);
        read(0, 55, 0, 0);
        nop(4);
        read(0, 55, 0, 0);
        nop(2);
        activate(5, 329);
        nop(2);
        read(0, 56, 0, 0);
        nop(4);
        read(0, 56, 0, 0);
        nop(4);
        read(0, 56, 0, 0);
        nop(4);
        read(0, 56, 0, 0);
        nop(4);
        read(5, 84, 0, 0);
        nop(4);
        read(5, 84, 0, 0);
        nop(4);
        read(5, 84, 0, 0);
        nop(4);
        read(5, 84, 0, 0);
        nop(4);
        read(5, 83, 0, 0);
        nop(4);
        read(0, 56, 0, 0);
        nop(2);
        precharge(5, 0);
        nop(2);
        read(0, 56, 0, 0);
        nop(4);
        read(0, 56, 0, 0);
        nop(4);
        read(0, 56, 0, 0);
        nop(2);
        activate(5, 503);
        nop(2);
        read(0, 57, 0, 0);
        nop(4);
        read(0, 57, 0, 0);
        nop(4);
        read(0, 57, 0, 0);
        nop(4);
        read(0, 57, 0, 0);
        nop(4);
        read(0, 57, 0, 0);
        nop(4);
        read(0, 57, 0, 0);
        nop(4);
        read(0, 57, 0, 0);
        nop(4);
        read(0, 57, 0, 0);
        nop(9);
        write(5, 85, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(5, 85, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(5, 85, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(5, 85, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(17);
        read(3, 108, 0, 0);
        nop(6);
        precharge(5, 0);
        nop(3);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(9);
        activate(5, 329);
        nop(8);
        read(3, 108, 0, 0);
        nop(4);
        read(5, 83, 0, 0);
        nop(4);
        read(5, 83, 0, 0);
        nop(4);
        read(5, 83, 0, 0);
        nop(4);
        read(5, 83, 0, 0);
        nop(4);
        read(5, 83, 0, 0);
        nop(4);
        read(5, 83, 0, 0);
        nop(4);
        read(5, 83, 0, 0);
        nop(4);
        read(5, 85, 0, 0);
        nop(4);
        read(5, 85, 0, 0);
        nop(4);
        read(5, 85, 0, 0);
        nop(4);
        read(5, 85, 0, 0);
        nop(4);
        read(5, 85, 0, 0);
        nop(4);
        read(5, 85, 0, 0);
        nop(4);
        read(5, 85, 0, 0);
        nop(4);
        read(5, 85, 0, 0);
        nop(9);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(17);
        read(3, 108, 0, 0);
        nop(9);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(17);
        read(3, 108, 0, 0);
        nop(9);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(202);
        precharge(2, 0);
        nop(12);
        activate(2, 369);
        nop(11);
        read(2, 52, 0, 0);
        nop(4);
        read(2, 52, 0, 0);
        nop(4);
        read(2, 52, 0, 0);
        nop(4);
        read(2, 52, 0, 0);
        nop(4);
        read(2, 52, 0, 0);
        nop(4);
        read(2, 52, 0, 0);
        nop(4);
        read(2, 52, 0, 0);
        nop(4);
        read(2, 52, 0, 0);
        nop(64);
        precharge(4, 0);
        nop(12);
        activate(4, 396);
        nop(11);
        read(4, 111, 0, 0);
        nop(4);
        read(4, 111, 0, 0);
        nop(4);
        read(4, 111, 0, 0);
        nop(4);
        read(4, 111, 0, 0);
        nop(4);
        read(4, 110, 0, 0);
        nop(6);
        precharge(4, 0);
        nop(3);
        precharge(7, 0);
        nop(9);
        activate(4, 396);
        nop(6);
        activate(7, 447);
        nop(5);
        read(4, 115, 0, 0);
        nop(4);
        read(4, 115, 0, 0);
        nop(4);
        read(4, 115, 0, 0);
        nop(2);
        precharge(5, 0);
        nop(2);
        read(4, 115, 0, 0);
        nop(4);
        read(4, 115, 0, 0);
        nop(4);
        read(7, 74, 0, 0);
        nop(2);
        precharge(4, 0);
        nop(1);
        activate(5, 396);
        nop(1);
        read(7, 74, 0, 0);
        nop(4);
        read(7, 74, 0, 0);
        nop(4);
        read(7, 74, 0, 0);
        nop(2);
        activate(4, 396);
        nop(2);
        read(5, 109, 0, 0);
        nop(4);
        read(5, 109, 0, 0);
        nop(4);
        read(7, 74, 0, 0);
        nop(4);
        read(7, 74, 0, 0);
        nop(4);
        read(4, 110, 0, 0);
        nop(4);
        read(4, 110, 0, 0);
        nop(4);
        read(4, 110, 0, 0);
        nop(4);
        read(4, 110, 0, 0);
        nop(4);
        read(4, 110, 0, 0);
        nop(4);
        read(5, 109, 0, 0);
        nop(2);
        precharge(4, 0);
        nop(2);
        read(7, 74, 0, 0);
        nop(4);
        read(5, 109, 0, 0);
        nop(4);
        read(7, 74, 0, 0);
        nop(2);
        activate(4, 396);
        nop(11);
        read(4, 115, 0, 0);
        nop(4);
        read(4, 115, 0, 0);
        nop(4);
        read(4, 115, 0, 0);
        nop(9);
        precharge(4, 0);
        nop(12);
        activate(4, 396);
        nop(11);
        read(4, 110, 0, 0);
        nop(4);
        read(4, 110, 0, 0);
        nop(4);
        read(4, 99, 0, 0);
        nop(4);
        read(4, 99, 0, 0);
        nop(4);
        read(4, 99, 0, 0);
        nop(6);
        precharge(4, 0);
        nop(12);
        activate(4, 394);
        nop(11);
        read(4, 87, 0, 0);
        nop(4);
        read(4, 87, 0, 0);
        nop(4);
        read(4, 87, 0, 0);
        nop(4);
        read(4, 87, 0, 0);
        nop(6);
        precharge(4, 0);
        nop(12);
        activate(4, 396);
        nop(11);
        read(4, 99, 0, 0);
        nop(4);
        read(4, 98, 0, 0);
        nop(4);
        read(4, 98, 0, 0);
        nop(4);
        read(4, 98, 0, 0);
        nop(4);
        read(4, 98, 0, 0);
        nop(6);
        precharge(4, 0);
        nop(12);
        activate(4, 394);
        nop(11);
        read(4, 90, 0, 0);
        nop(4);
        read(4, 90, 0, 0);
        nop(4);
        read(4, 90, 0, 0);
        nop(4);
        read(4, 90, 0, 0);
        nop(6);
        precharge(4, 0);
        nop(12);
        activate(4, 396);
        nop(11);
        read(4, 98, 0, 0);
        nop(4);
        read(4, 98, 0, 0);
        nop(4);
        read(4, 98, 0, 0);
        nop(4);
        read(4, 98, 0, 0);
        nop(2);
        precharge(0, 0);
        nop(2);
        read(4, 103, 0, 0);
        nop(6);
        precharge(4, 0);
        nop(4);
        activate(0, 17);
        nop(8);
        activate(4, 396);
        nop(3);
        read(0, 16, 0, 0);
        nop(4);
        read(0, 16, 0, 0);
        nop(4);
        read(0, 16, 0, 0);
        nop(4);
        read(0, 16, 0, 0);
        nop(4);
        read(0, 16, 0, 0);
        nop(4);
        read(0, 16, 0, 0);
        nop(4);
        read(3, 108, 0, 0);
        nop(4);
        read(4, 76, 0, 0);
        nop(4);
        read(4, 76, 0, 0);
        nop(4);
        read(4, 76, 0, 0);
        nop(4);
        read(0, 16, 0, 0);
        nop(4);
        read(0, 16, 0, 0);
        nop(4);
        read(4, 76, 0, 0);
        nop(4);
        read(4, 75, 0, 0);
        nop(6);
        precharge(4, 0);
        nop(3);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(9);
        activate(4, 396);
        nop(11);
        read(4, 103, 0, 0);
        nop(4);
        read(4, 103, 0, 0);
        nop(4);
        read(4, 103, 0, 0);
        nop(4);
        read(4, 103, 0, 0);
        nop(4);
        read(4, 103, 0, 0);
        nop(6);
        precharge(4, 0);
        nop(12);
        activate(4, 396);
        nop(11);
        read(4, 75, 0, 0);
        nop(4);
        read(4, 75, 0, 0);
        nop(4);
        read(3, 108, 0, 0);
        nop(4);
        read(4, 75, 0, 0);
        nop(6);
        precharge(4, 0);
        nop(3);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(9);
        activate(4, 396);
        nop(8);
        read(3, 108, 0, 0);
        nop(4);
        read(4, 103, 0, 0);
        nop(4);
        read(4, 103, 0, 0);
        nop(9);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(3);
        precharge(4, 0);
        nop(12);
        activate(4, 396);
        nop(11);
        read(4, 80, 0, 0);
        nop(4);
        read(4, 80, 0, 0);
        nop(4);
        read(4, 80, 0, 0);
        nop(4);
        read(4, 80, 0, 0);
        nop(4);
        read(4, 81, 0, 0);
        nop(6);
        precharge(4, 0);
        nop(12);
        activate(4, 408);
        nop(11);
        write(4, 80, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(4, 80, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(4, 80, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(4, 80, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(23);
        precharge(4, 0);
        nop(1);
        read(3, 108, 0, 0);
        nop(9);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(2);
        activate(4, 396);
        nop(2);
        precharge(0, 0);
        nop(12);
        activate(0, 321);
        nop(1);
        read(4, 81, 0, 0);
        nop(4);
        read(4, 81, 0, 0);
        nop(4);
        read(4, 81, 0, 0);
        nop(4);
        read(4, 81, 0, 0);
        nop(4);
        read(0, 58, 0, 0);
        nop(4);
        read(0, 58, 0, 0);
        nop(4);
        read(0, 58, 0, 0);
        nop(4);
        read(0, 58, 0, 0);
        nop(4);
        read(3, 108, 0, 0);
        nop(4);
        read(4, 81, 0, 0);
        nop(4);
        read(0, 58, 0, 0);
        nop(2);
        precharge(4, 0);
        nop(2);
        read(0, 58, 0, 0);
        nop(4);
        read(0, 58, 0, 0);
        nop(4);
        read(0, 58, 0, 0);
        nop(2);
        activate(4, 393);
        nop(7);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(17);
        read(4, 79, 0, 0);
        nop(4);
        read(4, 79, 0, 0);
        nop(4);
        read(4, 79, 0, 0);
        nop(4);
        read(4, 79, 0, 0);
        nop(6);
        precharge(4, 0);
        nop(12);
        activate(4, 396);
        nop(11);
        read(4, 81, 0, 0);
        nop(4);
        read(4, 81, 0, 0);
        nop(17);
        read(3, 108, 0, 0);
        nop(9);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(17);
        read(3, 108, 0, 0);
        nop(9);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(123);
        read(3, 108, 0, 0);
        nop(8);
        read(0, 60, 0, 0);
        nop(4);
        read(0, 60, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(2);
        read(0, 60, 0, 0);
        nop(4);
        read(0, 60, 0, 0);
        nop(1);
        precharge(1, 0);
        nop(5);
        activate(2, 461);
        nop(3);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        activate(1, 407);
        nop(13);
        read(1, 0, 0, 0);
        nop(4);
        read(1, 0, 0, 0);
        nop(4);
        read(2, 63, 0, 0);
        nop(4);
        read(1, 0, 0, 0);
        nop(4);
        read(1, 0, 0, 0);
        nop(4);
        read(1, 0, 0, 0);
        nop(4);
        read(1, 0, 0, 0);
        nop(2);
        precharge(0, 0);
        nop(2);
        read(1, 0, 0, 0);
        nop(4);
        read(1, 0, 0, 0);
        nop(4);
        read(2, 63, 0, 0);
        nop(2);
        activate(0, 1559);
        nop(2);
        read(1, 1, 0, 0);
        nop(4);
        read(1, 1, 0, 0);
        nop(4);
        read(1, 1, 0, 0);
        nop(4);
        read(0, 75, 0, 0);
        nop(2);
        precharge(5, 0);
        nop(2);
        read(1, 1, 0, 0);
        nop(4);
        read(2, 63, 0, 0);
        nop(4);
        read(0, 75, 0, 0);
        nop(2);
        activate(5, 363);
        nop(1);
        precharge(7, 0);
        nop(1);
        read(0, 75, 0, 0);
        nop(4);
        read(0, 75, 0, 0);
        nop(4);
        read(0, 75, 0, 0);
        nop(3);
        activate(7, 421);
        nop(1);
        read(2, 63, 0, 0);
        nop(4);
        read(0, 75, 0, 0);
        nop(4);
        read(0, 75, 0, 0);
        nop(4);
        read(7, 27, 0, 0);
        nop(4);
        read(7, 27, 0, 0);
        nop(4);
        read(7, 27, 0, 0);
        nop(4);
        read(0, 75, 0, 0);
        nop(4);
        read(1, 2, 0, 0);
        nop(4);
        read(7, 27, 0, 0);
        nop(4);
        read(7, 27, 0, 0);
        nop(4);
        read(1, 2, 0, 0);
        nop(2);
        precharge(7, 0);
        nop(2);
        read(1, 2, 0, 0);
        nop(4);
        read(1, 2, 0, 0);
        nop(4);
        read(1, 2, 0, 0);
        nop(2);
        activate(7, 930);
        nop(2);
        read(1, 2, 0, 0);
        nop(4);
        read(1, 2, 0, 0);
        nop(4);
        read(1, 2, 0, 0);
        nop(4);
        read(1, 3, 0, 0);
        nop(4);
        read(1, 3, 0, 0);
        nop(4);
        read(1, 3, 0, 0);
        nop(4);
        read(1, 3, 0, 0);
        nop(4);
        read(1, 3, 0, 0);
        nop(4);
        read(1, 3, 0, 0);
        nop(4);
        read(1, 3, 0, 0);
        nop(4);
        read(1, 3, 0, 0);
        nop(4);
        read(1, 4, 0, 0);
        nop(4);
        read(1, 4, 0, 0);
        nop(4);
        read(1, 4, 0, 0);
        nop(4);
        read(1, 4, 0, 0);
        nop(4);
        read(1, 5, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(2);
        read(1, 5, 0, 0);
        nop(4);
        read(1, 5, 0, 0);
        nop(4);
        read(1, 5, 0, 0);
        nop(2);
        activate(2, 407);
        nop(2);
        read(1, 6, 0, 0);
        nop(6);
        precharge(1, 0);
        nop(3);
        read(2, 78, 0, 0);
        nop(4);
        read(2, 78, 0, 0);
        nop(4);
        read(2, 78, 0, 0);
        nop(1);
        activate(1, 407);
        nop(3);
        read(2, 78, 0, 0);
        nop(8);
        read(1, 16, 0, 0);
        nop(4);
        read(1, 16, 0, 0);
        nop(4);
        read(1, 16, 0, 0);
        nop(4);
        read(1, 16, 0, 0);
        nop(4);
        read(1, 16, 0, 0);
        nop(6);
        precharge(1, 0);
        nop(3);
        write(5, 75, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(5, 75, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(7, 27, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(1);
        activate(1, 407);
        nop(3);
        write(5, 75, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(5, 75, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(7, 27, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(7, 27, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(7, 27, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(17);
        read(0, 76, 0, 0);
        nop(4);
        read(0, 76, 0, 0);
        nop(2);
        precharge(7, 0);
        nop(2);
        read(0, 76, 0, 0);
        nop(4);
        read(1, 6, 0, 0);
        nop(4);
        read(0, 76, 0, 0);
        nop(2);
        activate(7, 421);
        nop(2);
        read(0, 76, 0, 0);
        nop(4);
        read(0, 76, 0, 0);
        nop(4);
        read(0, 76, 0, 0);
        nop(4);
        read(7, 27, 0, 0);
        nop(4);
        read(0, 76, 0, 0);
        nop(4);
        read(1, 6, 0, 0);
        nop(4);
        read(7, 27, 0, 0);
        nop(2);
        precharge(5, 0);
        nop(2);
        read(7, 27, 0, 0);
        nop(4);
        read(1, 6, 0, 0);
        nop(4);
        read(1, 6, 0, 0);
        nop(2);
        activate(5, 441);
        nop(2);
        read(1, 6, 0, 0);
        nop(6);
        precharge(1, 0);
        nop(3);
        read(5, 76, 0, 0);
        nop(4);
        read(5, 76, 0, 0);
        nop(4);
        read(5, 76, 0, 0);
        nop(1);
        activate(1, 407);
        nop(3);
        read(5, 76, 0, 0);
        nop(6);
        precharge(5, 0);
        nop(2);
        read(1, 16, 0, 0);
        nop(4);
        read(1, 16, 0, 0);
        nop(4);
        read(1, 16, 0, 0);
        nop(2);
        activate(5, 363);
        nop(7);
        precharge(1, 0);
        nop(4);
        write(5, 76, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(5, 76, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        activate(1, 407);
        nop(1);
        write(5, 76, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(5, 76, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(17);
        read(1, 6, 0, 0);
        nop(4);
        read(1, 6, 0, 0);
        nop(2);
        precharge(5, 0);
        nop(2);
        read(1, 12, 0, 0);
        nop(4);
        read(1, 12, 0, 0);
        nop(4);
        read(1, 12, 0, 0);
        nop(2);
        activate(5, 441);
        nop(4);
        precharge(1, 0);
        nop(7);
        read(5, 76, 0, 0);
        nop(4);
        read(5, 76, 0, 0);
        nop(1);
        activate(1, 1419);
        nop(3);
        read(5, 76, 0, 0);
        nop(4);
        read(5, 76, 0, 0);
        nop(2);
        precharge(3, 0);
        nop(2);
        read(1, 73, 0, 0);
        nop(4);
        read(1, 73, 0, 0);
        nop(4);
        read(5, 75, 0, 0);
        nop(2);
        activate(3, 407);
        nop(2);
        read(5, 75, 0, 0);
        nop(4);
        read(5, 75, 0, 0);
        nop(4);
        read(1, 73, 0, 0);
        nop(4);
        read(1, 73, 0, 0);
        nop(4);
        read(1, 73, 0, 0);
        nop(4);
        read(3, 29, 0, 0);
        nop(2);
        precharge(1, 0);
        nop(2);
        read(3, 29, 0, 0);
        nop(4);
        read(5, 75, 0, 0);
        nop(4);
        read(3, 29, 0, 0);
        nop(2);
        activate(1, 407);
        nop(2);
        read(3, 29, 0, 0);
        nop(4);
        read(3, 31, 0, 0);
        nop(4);
        read(3, 31, 0, 0);
        nop(4);
        read(3, 31, 0, 0);
        nop(4);
        read(3, 31, 0, 0);
        nop(4);
        read(1, 12, 0, 0);
        nop(2);
        precharge(3, 0);
        nop(2);
        read(1, 13, 0, 0);
        nop(4);
        read(1, 13, 0, 0);
        nop(4);
        read(1, 13, 0, 0);
        nop(2);
        activate(3, 1585);
        nop(2);
        read(1, 13, 0, 0);
        nop(6);
        precharge(1, 0);
        nop(3);
        write(3, 31, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(3, 31, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(3, 31, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(1);
        activate(1, 1419);
        nop(3);
        write(3, 31, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(3, 31, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(3, 31, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(3, 31, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(3, 31, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(17);
        read(1, 73, 0, 0);
        nop(4);
        read(1, 73, 0, 0);
        nop(4);
        read(1, 73, 0, 0);
        nop(4);
        read(5, 66, 0, 0);
        nop(2);
        precharge(1, 0);
        nop(2);
        read(5, 66, 0, 0);
        nop(4);
        read(5, 66, 0, 0);
        nop(4);
        read(5, 66, 0, 0);
        nop(2);
        activate(1, 407);
        nop(4);
        precharge(5, 0);
        nop(7);
        read(1, 13, 0, 0);
        nop(4);
        read(1, 13, 0, 0);
        nop(1);
        activate(5, 452);
        nop(3);
        read(1, 13, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(2);
        read(1, 13, 0, 0);
        nop(4);
        read(5, 44, 0, 0);
        nop(4);
        read(1, 5, 0, 0);
        nop(2);
        activate(2, 499);
        nop(2);
        read(5, 44, 0, 0);
        nop(2);
        precharge(1, 0);
        nop(2);
        read(5, 44, 0, 0);
        nop(4);
        read(5, 44, 0, 0);
        nop(4);
        read(2, 67, 0, 0);
        nop(2);
        activate(1, 422);
        nop(2);
        read(2, 67, 0, 0);
        nop(4);
        read(2, 67, 0, 0);
        nop(4);
        read(2, 67, 0, 0);
        nop(4);
        read(1, 49, 0, 0);
        nop(4);
        read(2, 67, 0, 0);
        nop(2);
        precharge(3, 0);
        nop(2);
        read(1, 49, 0, 0);
        nop(4);
        read(1, 49, 0, 0);
        nop(4);
        read(1, 49, 0, 0);
        nop(2);
        activate(3, 407);
        nop(2);
        read(1, 49, 0, 0);
        nop(4);
        read(2, 67, 0, 0);
        nop(2);
        precharge(1, 0);
        nop(2);
        read(2, 67, 0, 0);
        nop(4);
        read(2, 67, 0, 0);
        nop(4);
        read(2, 66, 0, 0);
        nop(2);
        activate(1, 407);
        nop(2);
        read(3, 32, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(2);
        read(3, 32, 0, 0);
        nop(4);
        read(3, 32, 0, 0);
        nop(4);
        read(3, 32, 0, 0);
        nop(2);
        activate(2, 503);
        nop(2);
        read(1, 5, 0, 0);
        nop(4);
        read(1, 5, 0, 0);
        nop(4);
        read(1, 5, 0, 0);
        nop(4);
        read(1, 7, 0, 0);
        nop(4);
        read(1, 7, 0, 0);
        nop(4);
        read(2, 115, 0, 0);
        nop(2);
        precharge(1, 0);
        nop(2);
        read(2, 115, 0, 0);
        nop(4);
        read(2, 115, 0, 0);
        nop(4);
        read(2, 115, 0, 0);
        nop(2);
        activate(1, 422);
        nop(2);
        read(2, 115, 0, 0);
        nop(4);
        read(3, 32, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(1);
        precharge(4, 0);
        nop(1);
        read(3, 32, 0, 0);
        nop(4);
        read(1, 49, 0, 0);
        nop(4);
        read(1, 49, 0, 0);
        nop(2);
        activate(2, 499);
        nop(2);
        read(1, 49, 0, 0);
        nop(4);
        read(1, 50, 0, 0);
        nop(1);
        activate(4, 501);
        nop(3);
        read(3, 32, 0, 0);
        nop(4);
        read(1, 50, 0, 0);
        nop(4);
        read(2, 66, 0, 0);
        nop(2);
        precharge(1, 0);
        nop(2);
        read(2, 66, 0, 0);
        nop(4);
        read(2, 66, 0, 0);
        nop(4);
        read(3, 32, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(1);
        activate(1, 407);
        nop(1);
        read(4, 36, 0, 0);
        nop(2);
        precharge(3, 0);
        nop(2);
        read(4, 36, 0, 0);
        nop(4);
        read(4, 36, 0, 0);
        nop(2);
        activate(2, 503);
        nop(2);
        read(1, 7, 0, 0);
        nop(4);
        activate(3, 518);
        nop(1);
        read(4, 36, 0, 0);
        nop(4);
        read(4, 36, 0, 0);
        nop(4);
        read(1, 7, 0, 0);
        nop(4);
        read(1, 7, 0, 0);
        nop(4);
        read(1, 7, 0, 0);
        nop(4);
        read(1, 7, 0, 0);
        nop(4);
        read(2, 115, 0, 0);
        nop(2);
        precharge(1, 0);
        nop(2);
        read(3, 70, 0, 0);
        nop(4);
        read(4, 36, 0, 0);
        nop(4);
        read(2, 115, 0, 0);
        nop(2);
        activate(1, 422);
        nop(2);
        read(2, 115, 0, 0);
        nop(4);
        read(3, 70, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(2);
        read(3, 70, 0, 0);
        nop(4);
        read(3, 70, 0, 0);
        nop(4);
        read(4, 36, 0, 0);
        nop(2);
        activate(2, 735);
        nop(2);
        read(1, 50, 0, 0);
        nop(4);
        read(1, 50, 0, 0);
        nop(4);
        read(1, 50, 0, 0);
        nop(4);
        read(1, 50, 0, 0);
        nop(4);
        read(2, 101, 0, 0);
        nop(4);
        read(3, 70, 0, 0);
        nop(4);
        read(4, 36, 0, 0);
        nop(2);
        precharge(3, 0);
        nop(2);
        read(1, 50, 0, 0);
        nop(4);
        read(2, 101, 0, 0);
        nop(2);
        precharge(1, 0);
        nop(2);
        read(2, 101, 0, 0);
        nop(2);
        activate(3, 522);
        nop(2);
        read(2, 101, 0, 0);
        nop(4);
        read(2, 101, 0, 0);
        nop(2);
        activate(1, 407);
        nop(2);
        read(2, 101, 0, 0);
        nop(4);
        read(2, 101, 0, 0);
        nop(4);
        read(2, 101, 0, 0);
        nop(4);
        read(1, 7, 0, 0);
        nop(9);
        write(3, 70, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(3, 70, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(1);
        precharge(1, 0);
        nop(3);
        write(3, 70, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(3, 70, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(5);
        activate(1, 422);
        nop(12);
        read(1, 50, 0, 0);
        nop(6);
        precharge(3, 0);
        nop(10);
        precharge(1, 0);
        nop(2);
        activate(3, 518);
        nop(10);
        activate(1, 407);
        nop(1);
        read(3, 70, 0, 0);
        nop(10);
        read(1, 17, 0, 0);
        nop(1);
        precharge(7, 1);
        nop(1);
        precharge(0, 1);
        nop(1);
        precharge(2, 1);
        nop(1);
        precharge(4, 1);
        nop(1);
        precharge(5, 1);
        nop(1);
        precharge(6, 1);
        nop(1);
        precharge(3, 1);
        nop(10);
        precharge(1, 1);
        nop(101);
        activate(1, 407);
        nop(6);
        activate(3, 518);
        nop(5);
        read(1, 17, 0, 0);
        nop(4);
        read(1, 17, 0, 0);
        nop(4);
        read(3, 70, 0, 0);
        nop(4);
        read(1, 17, 0, 0);
        nop(4);
        read(1, 17, 0, 0);
        nop(4);
        read(1, 17, 0, 0);
        nop(4);
        read(1, 17, 0, 0);
        nop(4);
        read(1, 17, 0, 0);
        nop(4);
        read(1, 18, 0, 0);
        nop(4);
        read(3, 70, 0, 0);
        nop(4);
        read(1, 18, 0, 0);
        nop(2);
        precharge(3, 0);
        nop(2);
        read(1, 18, 0, 0);
        nop(4);
        read(1, 18, 0, 0);
        nop(4);
        read(1, 19, 0, 0);
        nop(2);
        activate(3, 521);
        nop(2);
        read(1, 19, 0, 0);
        nop(4);
        read(1, 19, 0, 0);
        nop(4);
        read(1, 19, 0, 0);
        nop(4);
        read(1, 19, 0, 0);
        nop(4);
        read(1, 19, 0, 0);
        nop(4);
        read(1, 19, 0, 0);
        nop(4);
        read(1, 19, 0, 0);
        nop(4);
        read(1, 20, 0, 0);
        nop(4);
        read(1, 20, 0, 0);
        nop(4);
        read(3, 43, 0, 0);
        nop(4);
        read(3, 43, 0, 0);
        nop(4);
        read(1, 20, 0, 0);
        nop(4);
        read(1, 20, 0, 0);
        nop(4);
        read(1, 20, 0, 0);
        nop(4);
        read(1, 20, 0, 0);
        nop(4);
        read(1, 20, 0, 0);
        nop(4);
        read(1, 20, 0, 0);
        nop(4);
        read(3, 43, 0, 0);
        nop(4);
        read(3, 43, 0, 0);
        nop(4);
        read(1, 22, 0, 0);
        nop(4);
        read(1, 22, 0, 0);
        nop(4);
        read(1, 22, 0, 0);
        nop(4);
        read(1, 22, 0, 0);
        nop(4);
        read(3, 42, 0, 0);
        nop(2);
        precharge(1, 0);
        nop(2);
        read(3, 42, 0, 0);
        nop(4);
        read(3, 42, 0, 0);
        nop(4);
        read(3, 42, 0, 0);
        nop(2);
        activate(1, 407);
        nop(11);
        read(1, 35, 0, 0);
        nop(4);
        read(1, 35, 0, 0);
        nop(4);
        read(1, 35, 0, 0);
        nop(4);
        read(1, 35, 0, 0);
        nop(4);
        read(1, 36, 0, 0);
        nop(6);
        precharge(1, 0);
        nop(12);
        activate(1, 407);
        nop(11);
        read(1, 22, 0, 0);
        nop(4);
        read(1, 22, 0, 0);
        nop(4);
        read(1, 22, 0, 0);
        nop(2);
        activate(0, 321);
        nop(2);
        read(1, 22, 0, 0);
        nop(4);
        read(1, 21, 0, 0);
        nop(5);
        read(0, 61, 0, 0);
        nop(1);
        precharge(1, 0);
        nop(3);
        read(0, 61, 0, 0);
        nop(4);
        read(0, 61, 0, 0);
        nop(4);
        read(0, 61, 0, 0);
        nop(1);
        activate(1, 407);
        nop(3);
        read(0, 61, 0, 0);
        nop(4);
        read(0, 61, 0, 0);
        nop(4);
        read(0, 61, 0, 0);
        nop(4);
        read(0, 61, 0, 0);
        nop(4);
        read(1, 36, 0, 0);
        nop(4);
        read(1, 36, 0, 0);
        nop(4);
        read(1, 36, 0, 0);
        nop(4);
        read(1, 36, 0, 0);
        nop(4);
        read(1, 36, 0, 0);
        nop(6);
        precharge(1, 0);
        nop(12);
        activate(1, 407);
        nop(11);
        read(1, 21, 0, 0);
        nop(2);
        activate(7, 459);
        nop(2);
        read(1, 21, 0, 0);
        nop(4);
        read(1, 21, 0, 0);
        nop(4);
        read(1, 23, 0, 0);
        nop(4);
        read(1, 23, 0, 0);
        nop(4);
        read(7, 28, 0, 0);
        nop(2);
        precharge(1, 0);
        nop(2);
        read(7, 28, 0, 0);
        nop(4);
        read(7, 28, 0, 0);
        nop(4);
        read(7, 28, 0, 0);
        nop(2);
        activate(1, 407);
        nop(2);
        read(7, 28, 0, 0);
        nop(6);
        precharge(7, 0);
        nop(3);
        read(1, 36, 0, 0);
        nop(4);
        read(1, 36, 0, 0);
        nop(5);
        activate(7, 450);
        nop(8);
        precharge(1, 0);
        nop(3);
        write(7, 28, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(7, 28, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(7, 28, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(1);
        activate(1, 407);
        nop(3);
        write(7, 28, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(17);
        read(1, 23, 0, 0);
        nop(4);
        read(1, 23, 0, 0);
        nop(2);
        precharge(7, 0);
        nop(2);
        read(1, 26, 0, 0);
        nop(4);
        read(1, 26, 0, 0);
        nop(2);
        activate(4, 317);
        nop(2);
        read(1, 26, 0, 0);
        nop(4);
        activate(7, 459);
        nop(2);
        precharge(1, 0);
        nop(3);
        read(4, 70, 0, 0);
        nop(4);
        read(4, 70, 0, 0);
        nop(4);
        read(7, 28, 0, 0);
        nop(1);
        activate(1, 1587);
        nop(3);
        read(4, 70, 0, 0);
        nop(4);
        read(4, 70, 0, 0);
        nop(4);
        read(4, 70, 0, 0);
        nop(4);
        read(4, 70, 0, 0);
        nop(4);
        read(4, 70, 0, 0);
        nop(4);
        read(7, 28, 0, 0);
        nop(4);
        read(7, 28, 0, 0);
        nop(4);
        read(7, 29, 0, 0);
        nop(4);
        read(1, 4, 0, 0);
        nop(4);
        read(1, 4, 0, 0);
        nop(4);
        read(4, 70, 0, 0);
        nop(4);
        read(7, 29, 0, 0);
        nop(4);
        read(1, 4, 0, 0);
        nop(2);
        precharge(7, 0);
        nop(2);
        read(1, 4, 0, 0);
        nop(4);
        read(1, 5, 0, 0);
        nop(6);
        precharge(1, 0);
        nop(1);
        activate(7, 459);
        nop(11);
        read(7, 40, 0, 0);
        nop(1);
        activate(1, 407);
        nop(3);
        read(7, 40, 0, 0);
        nop(4);
        read(7, 40, 0, 0);
        nop(4);
        read(7, 40, 0, 0);
        nop(4);
        read(7, 41, 0, 0);
        nop(4);
        read(1, 26, 0, 0);
        nop(2);
        precharge(7, 0);
        nop(2);
        read(1, 26, 0, 0);
        nop(4);
        read(1, 26, 0, 0);
        nop(4);
        read(1, 26, 0, 0);
        nop(2);
        activate(7, 459);
        nop(2);
        read(1, 26, 0, 0);
        nop(6);
        precharge(1, 0);
        nop(3);
        read(7, 29, 0, 0);
        nop(4);
        read(7, 29, 0, 0);
        nop(4);
        read(7, 29, 0, 0);
        nop(1);
        activate(1, 1587);
        nop(3);
        read(7, 29, 0, 0);
        nop(4);
        read(7, 29, 0, 0);
        nop(4);
        read(1, 5, 0, 0);
        nop(2);
        precharge(7, 0);
        nop(2);
        read(1, 5, 0, 0);
        nop(2);
        activate(5, 1581);
        nop(2);
        read(1, 5, 0, 0);
        nop(6);
        activate(7, 459);
        nop(3);
        read(5, 126, 0, 0);
        nop(1);
        precharge(1, 0);
        nop(3);
        read(5, 126, 0, 0);
        nop(4);
        read(7, 41, 0, 0);
        nop(4);
        read(5, 126, 0, 0);
        nop(1);
        activate(1, 407);
        nop(3);
        read(5, 126, 0, 0);
        nop(4);
        read(5, 126, 0, 0);
        nop(4);
        read(5, 126, 0, 0);
        nop(4);
        read(7, 41, 0, 0);
        nop(2);
        precharge(5, 0);
        nop(2);
        read(7, 41, 0, 0);
        nop(4);
        read(1, 30, 0, 0);
        nop(4);
        read(1, 30, 0, 0);
        nop(2);
        activate(5, 928);
        nop(2);
        read(7, 41, 0, 0);
        nop(4);
        read(7, 41, 0, 0);
        nop(4);
        read(1, 30, 0, 0);
        nop(2);
        precharge(7, 0);
        nop(2);
        read(1, 30, 0, 0);
        nop(4);
        read(1, 30, 0, 0);
        nop(4);
        read(1, 30, 0, 0);
        nop(2);
        activate(7, 459);
        nop(2);
        read(1, 30, 0, 0);
        nop(4);
        read(1, 30, 0, 0);
        nop(5);
        read(7, 29, 0, 0);
        nop(9);
        write(5, 126, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(5, 126, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(5, 126, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(1);
        precharge(7, 0);
        nop(3);
        write(5, 126, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(9);
        activate(7, 459);
        nop(11);
        read(7, 41, 0, 0);
        nop(3);
        precharge(5, 0);
        nop(1);
        read(7, 41, 0, 0);
        nop(4);
        read(7, 42, 0, 0);
        nop(4);
        read(7, 42, 0, 0);
        nop(3);
        activate(5, 1581);
        nop(1);
        read(7, 42, 0, 0);
        nop(6);
        precharge(7, 0);
        nop(4);
        read(5, 126, 0, 0);
        nop(4);
        read(5, 126, 0, 0);
        nop(4);
        activate(7, 425);
        nop(1);
        read(5, 127, 0, 0);
        nop(4);
        read(5, 127, 0, 0);
        nop(4);
        read(5, 127, 0, 0);
        nop(4);
        read(5, 127, 0, 0);
        nop(4);
        read(5, 127, 0, 0);
        nop(4);
        read(5, 127, 0, 0);
        nop(4);
        read(5, 127, 0, 0);
        nop(4);
        read(5, 127, 0, 0);
        nop(9);
        write(7, 41, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(7, 41, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(7, 41, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(7, 41, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(23);
        precharge(7, 0);
        nop(12);
        activate(7, 459);
        nop(11);
        read(7, 42, 0, 0);
        nop(4);
        read(7, 42, 0, 0);
        nop(4);
        read(7, 42, 0, 0);
        nop(4);
        read(7, 42, 0, 0);
        nop(4);
        read(7, 42, 0, 0);
        nop(6);
        precharge(7, 0);
        nop(12);
        activate(7, 449);
        nop(11);
        write(7, 42, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(7, 42, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(7, 42, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(7, 42, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(23);
        precharge(7, 0);
        nop(12);
        activate(7, 421);
        nop(11);
        read(7, 0, 0, 0);
        nop(4);
        read(7, 0, 0, 0);
        nop(4);
        read(7, 0, 0, 0);
        nop(4);
        read(7, 0, 0, 0);
        nop(4);
        read(7, 0, 0, 0);
        nop(6);
        precharge(7, 0);
        nop(12);
        activate(7, 459);
        nop(11);
        read(7, 52, 0, 0);
        nop(4);
        read(7, 52, 0, 0);
        nop(4);
        read(7, 52, 0, 0);
        nop(4);
        read(7, 52, 0, 0);
        nop(4);
        read(7, 53, 0, 0);
        nop(6);
        precharge(7, 0);
        nop(12);
        activate(7, 421);
        nop(11);
        read(7, 0, 0, 0);
        nop(4);
        read(7, 0, 0, 0);
        nop(4);
        read(7, 0, 0, 0);
        nop(4);
        read(7, 2, 0, 0);
        nop(4);
        read(7, 2, 0, 0);
        nop(6);
        precharge(7, 0);
        nop(12);
        activate(7, 459);
        nop(11);
        read(7, 53, 0, 0);
        nop(4);
        read(7, 53, 0, 0);
        nop(4);
        read(7, 53, 0, 0);
        nop(4);
        read(7, 53, 0, 0);
        nop(4);
        read(7, 53, 0, 0);
        nop(6);
        precharge(7, 0);
        nop(12);
        activate(7, 421);
        nop(11);
        read(7, 2, 0, 0);
        nop(4);
        read(7, 2, 0, 0);
        nop(4);
        read(7, 3, 0, 0);
        nop(4);
        read(7, 3, 0, 0);
        nop(4);
        read(7, 3, 0, 0);
        nop(6);
        precharge(7, 0);
        nop(12);
        activate(7, 459);
        nop(11);
        read(7, 53, 0, 0);
        nop(4);
        read(7, 53, 0, 0);
        nop(4);
        read(7, 54, 0, 0);
        nop(4);
        read(7, 54, 0, 0);
        nop(4);
        read(7, 54, 0, 0);
        nop(6);
        precharge(7, 0);
        nop(12);
        activate(7, 421);
        nop(11);
        read(7, 3, 0, 0);
        nop(4);
        read(7, 3, 0, 0);
        nop(4);
        read(7, 3, 0, 0);
        nop(4);
        read(7, 3, 0, 0);
        nop(4);
        read(7, 3, 0, 0);
        nop(6);
        precharge(7, 0);
        nop(12);
        activate(7, 459);
        nop(11);
        read(7, 12, 0, 0);
        nop(4);
        read(7, 12, 0, 0);
        nop(4);
        read(7, 12, 0, 0);
        nop(4);
        read(7, 12, 0, 0);
        nop(6);
        precharge(7, 0);
        nop(12);
        activate(7, 459);
        nop(11);
        read(7, 54, 0, 0);
        nop(4);
        read(7, 55, 0, 0);
        nop(4);
        read(7, 55, 0, 0);
        nop(4);
        read(7, 55, 0, 0);
        nop(4);
        read(7, 55, 0, 0);
        nop(4);
        read(0, 62, 0, 0);
        nop(2);
        precharge(7, 0);
        nop(2);
        read(0, 62, 0, 0);
        nop(4);
        read(0, 62, 0, 0);
        nop(2);
        activate(2, 461);
        nop(2);
        read(0, 62, 0, 0);
        nop(4);
        activate(7, 510);
        nop(5);
        read(2, 83, 0, 0);
        nop(4);
        read(2, 83, 0, 0);
        nop(4);
        read(2, 83, 0, 0);
        nop(4);
        read(2, 83, 0, 0);
        nop(4);
        read(2, 83, 0, 0);
        nop(4);
        read(2, 83, 0, 0);
        nop(4);
        read(2, 83, 0, 0);
        nop(4);
        read(2, 83, 0, 0);
        nop(4);
        read(2, 89, 0, 0);
        nop(4);
        read(2, 89, 0, 0);
        nop(4);
        read(2, 89, 0, 0);
        nop(4);
        read(2, 89, 0, 0);
        nop(4);
        read(2, 90, 0, 0);
        nop(4);
        read(2, 90, 0, 0);
        nop(4);
        read(2, 90, 0, 0);
        nop(4);
        read(2, 90, 0, 0);
        nop(4);
        read(2, 91, 0, 0);
        nop(4);
        read(2, 91, 0, 0);
        nop(4);
        read(2, 91, 0, 0);
        nop(4);
        read(2, 91, 0, 0);
        nop(4);
        read(2, 91, 0, 0);
        nop(4);
        read(2, 91, 0, 0);
        nop(4);
        read(2, 91, 0, 0);
        nop(4);
        read(2, 91, 0, 0);
        nop(4);
        read(2, 93, 0, 0);
        nop(4);
        read(2, 93, 0, 0);
        nop(4);
        read(2, 93, 0, 0);
        nop(4);
        read(2, 93, 0, 0);
        nop(4);
        read(2, 93, 0, 0);
        nop(4);
        read(2, 93, 0, 0);
        nop(4);
        read(2, 93, 0, 0);
        nop(2);
        precharge(3, 0);
        nop(2);
        read(2, 93, 0, 0);
        nop(9);
        write(7, 55, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(1);
        activate(3, 2026);
        nop(3);
        write(7, 55, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(7, 55, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(7, 55, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(7, 55, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(17);
        read(3, 108, 0, 0);
        nop(6);
        precharge(7, 0);
        nop(3);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(9);
        activate(7, 459);
        nop(8);
        read(3, 108, 0, 0);
        nop(4);
        read(7, 55, 0, 0);
        nop(4);
        read(7, 55, 0, 0);
        nop(4);
        read(7, 55, 0, 0);
        nop(4);
        read(7, 55, 0, 0);
        nop(4);
        read(7, 56, 0, 0);
        nop(6);
        precharge(7, 0);
        nop(3);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(9);
        activate(7, 510);
        nop(8);
        read(3, 108, 0, 0);
        nop(2);
        precharge(4, 0);
        nop(7);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(7, 55, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(1);
        activate(4, 482);
        nop(3);
        write(7, 55, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(7, 55, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(17);
        read(3, 108, 0, 0);
        nop(4);
        read(4, 73, 0, 0);
        nop(2);
        precharge(7, 0);
        nop(2);
        read(4, 73, 0, 0);
        nop(2);
        precharge(5, 0);
        nop(2);
        read(4, 73, 0, 0);
        nop(4);
        read(4, 73, 0, 0);
        nop(2);
        activate(7, 459);
        nop(2);
        read(4, 73, 0, 0);
        nop(4);
        read(4, 73, 0, 0);
        nop(1);
        activate(5, 1831);
        nop(3);
        read(4, 73, 0, 0);
        nop(4);
        read(4, 73, 0, 0);
        nop(4);
        read(5, 6, 0, 0);
        nop(4);
        read(7, 56, 0, 0);
        nop(4);
        read(7, 56, 0, 0);
        nop(4);
        read(5, 6, 0, 0);
        nop(4);
        read(5, 6, 0, 0);
        nop(4);
        read(5, 6, 0, 0);
        nop(4);
        read(7, 56, 0, 0);
        nop(2);
        precharge(5, 0);
        nop(2);
        read(7, 57, 0, 0);
        nop(4);
        read(7, 57, 0, 0);
        nop(6);
        precharge(7, 0);
        nop(1);
        activate(5, 422);
        nop(2);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(9);
        activate(7, 930);
        nop(8);
        read(3, 108, 0, 0);
        nop(4);
        read(5, 65, 0, 0);
        nop(4);
        read(5, 65, 0, 0);
        nop(4);
        read(5, 65, 0, 0);
        nop(2);
        precharge(4, 0);
        nop(2);
        read(5, 65, 0, 0);
        nop(4);
        read(5, 65, 0, 0);
        nop(4);
        read(5, 65, 0, 0);
        nop(2);
        activate(4, 386);
        nop(1);
        precharge(1, 0);
        nop(1);
        read(5, 65, 0, 0);
        nop(4);
        read(5, 65, 0, 0);
        nop(5);
        read(4, 37, 0, 0);
        nop(2);
        activate(1, 407);
        nop(2);
        read(4, 37, 0, 0);
        nop(4);
        read(4, 37, 0, 0);
        nop(4);
        read(4, 37, 0, 0);
        nop(4);
        read(4, 37, 0, 0);
        nop(4);
        read(1, 39, 0, 0);
        nop(4);
        read(1, 39, 0, 0);
        nop(4);
        read(1, 39, 0, 0);
        nop(4);
        read(1, 39, 0, 0);
        nop(4);
        read(4, 37, 0, 0);
        nop(2);
        precharge(1, 0);
        nop(2);
        read(4, 37, 0, 0);
        nop(4);
        read(4, 37, 0, 0);
        nop(6);
        activate(1, 405);
        nop(3);
        write(7, 56, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(7, 56, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(2);
        precharge(0, 0);
        nop(2);
        write(7, 56, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(7, 56, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(6);
        activate(0, 1558);
        nop(11);
        read(0, 111, 0, 0);
        nop(4);
        read(0, 111, 0, 0);
        nop(2);
        precharge(7, 0);
        nop(2);
        read(0, 111, 0, 0);
        nop(4);
        read(1, 50, 0, 0);
        nop(4);
        read(3, 108, 0, 0);
        nop(2);
        activate(7, 459);
        nop(2);
        read(0, 111, 0, 0);
        nop(4);
        read(0, 111, 0, 0);
        nop(4);
        read(0, 111, 0, 0);
        nop(4);
        read(7, 57, 0, 0);
        nop(4);
        read(0, 111, 0, 0);
        nop(4);
        read(1, 50, 0, 0);
        nop(4);
        read(7, 57, 0, 0);
        nop(4);
        read(7, 57, 0, 0);
        nop(4);
        read(7, 57, 0, 0);
        nop(4);
        read(7, 57, 0, 0);
        nop(4);
        read(0, 111, 0, 0);
        nop(2);
        precharge(7, 0);
        nop(2);
        read(1, 50, 0, 0);
        nop(4);
        read(1, 50, 0, 0);
        nop(4);
        read(1, 50, 0, 0);
        nop(2);
        activate(7, 421);
        nop(4);
        precharge(1, 0);
        nop(3);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(9);
        activate(1, 407);
        nop(8);
        read(7, 97, 0, 0);
        nop(4);
        read(1, 37, 0, 0);
        nop(4);
        read(1, 37, 0, 0);
        nop(4);
        read(3, 108, 0, 0);
        nop(4);
        read(4, 35, 0, 0);
        nop(4);
        read(4, 35, 0, 0);
        nop(4);
        read(7, 97, 0, 0);
        nop(4);
        read(7, 97, 0, 0);
        nop(4);
        read(7, 97, 0, 0);
        nop(4);
        read(1, 37, 0, 0);
        nop(4);
        read(1, 37, 0, 0);
        nop(4);
        read(4, 35, 0, 0);
        nop(4);
        read(4, 35, 0, 0);
        nop(4);
        read(7, 97, 0, 0);
        nop(4);
        read(1, 37, 0, 0);
        nop(2);
        precharge(7, 0);
        nop(4);
        precharge(1, 0);
        nop(3);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(5);
        activate(7, 459);
        nop(6);
        activate(1, 405);
        nop(6);
        read(3, 108, 0, 0);
        nop(4);
        read(7, 57, 0, 0);
        nop(4);
        read(7, 58, 0, 0);
        nop(4);
        read(7, 58, 0, 0);
        nop(4);
        read(7, 58, 0, 0);
        nop(4);
        read(1, 50, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(2);
        read(7, 58, 0, 0);
        nop(4);
        read(1, 50, 0, 0);
        nop(2);
        precharge(7, 0);
        nop(2);
        read(1, 50, 0, 0);
        nop(2);
        activate(2, 423);
        nop(2);
        read(1, 51, 0, 0);
        nop(4);
        read(1, 51, 0, 0);
        nop(2);
        activate(7, 421);
        nop(3);
        read(2, 56, 0, 0);
        nop(1);
        precharge(1, 0);
        nop(3);
        read(2, 56, 0, 0);
        nop(4);
        read(7, 97, 0, 0);
        nop(4);
        read(7, 97, 0, 0);
        nop(1);
        activate(1, 407);
        nop(3);
        read(2, 56, 0, 0);
        nop(4);
        read(2, 56, 0, 0);
        nop(4);
        read(2, 56, 0, 0);
        nop(4);
        read(7, 97, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(2);
        read(1, 37, 0, 0);
        nop(4);
        read(1, 37, 0, 0);
        nop(4);
        read(1, 37, 0, 0);
        nop(2);
        activate(2, 930);
        nop(2);
        read(1, 38, 0, 0);
        nop(4);
        read(1, 38, 0, 0);
        nop(6);
        precharge(1, 0);
        nop(3);
        write(2, 56, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(2, 56, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(2, 56, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(1);
        activate(1, 405);
        nop(3);
        write(2, 56, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(17);
        read(1, 51, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(2);
        read(1, 51, 0, 0);
        nop(4);
        read(1, 51, 0, 0);
        nop(4);
        read(1, 51, 0, 0);
        nop(2);
        activate(2, 423);
        nop(2);
        read(1, 51, 0, 0);
        nop(6);
        precharge(1, 0);
        nop(3);
        read(2, 56, 0, 0);
        nop(4);
        read(2, 56, 0, 0);
        nop(4);
        read(2, 56, 0, 0);
        nop(1);
        activate(1, 407);
        nop(3);
        read(2, 61, 0, 0);
        nop(4);
        read(2, 61, 0, 0);
        nop(4);
        read(1, 38, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(2);
        read(1, 38, 0, 0);
        nop(4);
        read(1, 38, 0, 0);
        nop(4);
        read(1, 38, 0, 0);
        nop(2);
        activate(2, 265);
        nop(2);
        read(1, 38, 0, 0);
        nop(6);
        precharge(1, 0);
        nop(3);
        read(2, 37, 0, 0);
        nop(4);
        read(2, 37, 0, 0);
        nop(4);
        read(2, 37, 0, 0);
        nop(1);
        activate(1, 405);
        nop(3);
        read(2, 37, 0, 0);
        nop(4);
        read(2, 37, 0, 0);
        nop(4);
        read(1, 51, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(12);
        activate(2, 423);
        nop(3);
        precharge(1, 0);
        nop(8);
        read(2, 61, 0, 0);
        nop(4);
        activate(1, 407);
        nop(1);
        read(2, 61, 0, 0);
        nop(4);
        read(2, 62, 0, 0);
        nop(4);
        read(2, 62, 0, 0);
        nop(4);
        read(1, 38, 0, 0);
        nop(4);
        read(1, 40, 0, 0);
        nop(4);
        read(1, 40, 0, 0);
        nop(4);
        read(2, 62, 0, 0);
        nop(4);
        read(1, 40, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(2);
        read(1, 40, 0, 0);
        nop(6);
        precharge(1, 0);
        nop(4);
        activate(2, 265);
        nop(8);
        activate(1, 407);
        nop(3);
        read(2, 37, 0, 0);
        nop(4);
        read(2, 37, 0, 0);
        nop(4);
        read(1, 64, 0, 0);
        nop(4);
        read(1, 64, 0, 0);
        nop(4);
        read(1, 64, 0, 0);
        nop(4);
        read(1, 64, 0, 0);
        nop(4);
        read(1, 64, 0, 0);
        nop(4);
        read(2, 37, 0, 0);
        nop(2);
        precharge(1, 0);
        nop(4);
        precharge(2, 0);
        nop(8);
        activate(1, 407);
        nop(6);
        activate(2, 511);
        nop(5);
        read(1, 40, 0, 0);
        nop(4);
        read(1, 40, 0, 0);
        nop(4);
        read(1, 40, 0, 0);
        nop(4);
        read(1, 40, 0, 0);
        nop(4);
        read(1, 41, 0, 0);
        nop(6);
        precharge(1, 0);
        nop(3);
        write(2, 61, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(2, 61, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(2, 61, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(1);
        activate(1, 407);
        nop(3);
        write(2, 61, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(17);
        read(1, 64, 0, 0);
        nop(4);
        read(1, 64, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(2);
        read(1, 64, 0, 0);
        nop(4);
        read(1, 65, 0, 0);
        nop(4);
        read(1, 65, 0, 0);
        nop(2);
        activate(2, 423);
        nop(4);
        precharge(1, 0);
        nop(7);
        read(2, 62, 0, 0);
        nop(4);
        read(2, 62, 0, 0);
        nop(1);
        activate(1, 407);
        nop(3);
        read(2, 62, 0, 0);
        nop(4);
        read(2, 62, 0, 0);
        nop(4);
        read(1, 41, 0, 0);
        nop(4);
        read(1, 41, 0, 0);
        nop(4);
        read(1, 41, 0, 0);
        nop(4);
        read(1, 41, 0, 0);
        nop(4);
        read(1, 41, 0, 0);
        nop(4);
        read(2, 62, 0, 0);
        nop(2);
        precharge(1, 0);
        nop(4);
        precharge(2, 0);
        nop(8);
        activate(1, 407);
        nop(6);
        activate(2, 500);
        nop(5);
        read(1, 65, 0, 0);
        nop(4);
        read(1, 65, 0, 0);
        nop(9);
        write(2, 63, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(2);
        precharge(7, 0);
        nop(2);
        precharge(1, 0);
        nop(1);
        write(2, 63, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(2, 63, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(2, 63, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(1);
        activate(7, 459);
        nop(6);
        activate(1, 407);
        nop(10);
        read(7, 0, 0, 0);
        nop(4);
        read(7, 0, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(2);
        read(7, 0, 0, 0);
        nop(4);
        read(7, 0, 0, 0);
        nop(4);
        read(7, 0, 0, 0);
        nop(2);
        activate(2, 423);
        nop(2);
        read(1, 41, 0, 0);
        nop(4);
        read(1, 41, 0, 0);
        nop(4);
        read(7, 0, 0, 0);
        nop(4);
        read(7, 0, 0, 0);
        nop(4);
        read(7, 0, 0, 0);
        nop(4);
        read(7, 1, 0, 0);
        nop(4);
        read(7, 1, 0, 0);
        nop(4);
        read(7, 1, 0, 0);
        nop(2);
        precharge(4, 0);
        nop(2);
        read(2, 51, 0, 0);
        nop(4);
        read(2, 51, 0, 0);
        nop(4);
        read(7, 1, 0, 0);
        nop(2);
        activate(4, 394);
        nop(2);
        read(7, 1, 0, 0);
        nop(4);
        read(7, 1, 0, 0);
        nop(4);
        read(7, 1, 0, 0);
        nop(4);
        read(2, 51, 0, 0);
        nop(4);
        read(2, 51, 0, 0);
        nop(4);
        read(2, 51, 0, 0);
        nop(4);
        read(4, 89, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(2);
        read(7, 1, 0, 0);
        nop(4);
        read(4, 89, 0, 0);
        nop(2);
        activate(6, 406);
        nop(2);
        read(4, 89, 0, 0);
        nop(4);
        activate(2, 405);
        nop(1);
        read(4, 89, 0, 0);
        nop(4);
        read(6, 33, 0, 0);
        nop(4);
        read(6, 33, 0, 0);
        nop(4);
        read(6, 33, 0, 0);
        nop(4);
        read(6, 33, 0, 0);
        nop(4);
        read(7, 4, 0, 0);
        nop(4);
        read(2, 10, 0, 0);
        nop(4);
        read(2, 10, 0, 0);
        nop(4);
        read(2, 10, 0, 0);
        nop(4);
        read(7, 4, 0, 0);
        nop(4);
        read(7, 4, 0, 0);
        nop(4);
        read(7, 4, 0, 0);
        nop(4);
        read(7, 2, 0, 0);
        nop(4);
        read(7, 2, 0, 0);
        nop(4);
        read(2, 10, 0, 0);
        nop(4);
        read(2, 15, 0, 0);
        nop(4);
        read(7, 2, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(4);
        precharge(7, 0);
        nop(8);
        activate(2, 423);
        nop(6);
        activate(7, 510);
        nop(5);
        read(2, 51, 0, 0);
        nop(4);
        read(2, 51, 0, 0);
        nop(4);
        read(2, 51, 0, 0);
        nop(4);
        read(2, 52, 0, 0);
        nop(4);
        read(2, 52, 0, 0);
        nop(6);
        precharge(2, 0);
        nop(3);
        write(7, 2, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(7, 2, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(7, 2, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(1);
        activate(2, 405);
        nop(3);
        write(7, 2, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(7, 2, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(17);
        read(1, 42, 0, 0);
        nop(4);
        read(1, 42, 0, 0);
        nop(2);
        precharge(7, 0);
        nop(2);
        read(1, 42, 0, 0);
        nop(4);
        read(1, 42, 0, 0);
        nop(4);
        read(1, 42, 0, 0);
        nop(2);
        activate(7, 459);
        nop(2);
        read(2, 15, 0, 0);
        nop(4);
        read(3, 108, 0, 0);
        nop(4);
        read(5, 66, 0, 0);
        nop(4);
        read(5, 66, 0, 0);
        nop(4);
        read(7, 2, 0, 0);
        nop(4);
        read(7, 2, 0, 0);
        nop(4);
        read(1, 42, 0, 0);
        nop(4);
        read(1, 42, 0, 0);
        nop(4);
        read(2, 15, 0, 0);
        nop(4);
        read(5, 66, 0, 0);
        nop(4);
        read(5, 66, 0, 0);
        nop(4);
        read(5, 67, 0, 0);
        nop(4);
        read(7, 2, 0, 0);
        nop(4);
        read(7, 2, 0, 0);
        nop(4);
        read(1, 42, 0, 0);
        nop(4);
        read(2, 15, 0, 0);
        nop(2);
        precharge(1, 0);
        nop(2);
        read(5, 67, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(2);
        read(5, 67, 0, 0);
        nop(4);
        read(7, 2, 0, 0);
        nop(2);
        activate(1, 265);
        nop(2);
        read(5, 67, 0, 0);
        nop(2);
        precharge(7, 0);
        nop(2);
        activate(2, 423);
        nop(1);
        read(5, 67, 0, 0);
        nop(4);
        read(5, 67, 0, 0);
        nop(4);
        read(5, 67, 0, 0);
        nop(1);
        activate(7, 510);
        nop(3);
        read(1, 70, 0, 0);
        nop(4);
        read(1, 70, 0, 0);
        nop(4);
        read(1, 70, 0, 0);
        nop(4);
        read(2, 52, 0, 0);
        nop(4);
        read(5, 67, 0, 0);
        nop(4);
        read(5, 68, 0, 0);
        nop(4);
        read(5, 68, 0, 0);
        nop(4);
        read(1, 70, 0, 0);
        nop(4);
        read(1, 71, 0, 0);
        nop(4);
        read(1, 71, 0, 0);
        nop(4);
        read(1, 71, 0, 0);
        nop(4);
        read(2, 52, 0, 0);
        nop(4);
        read(5, 68, 0, 0);
        nop(4);
        read(5, 68, 0, 0);
        nop(4);
        read(5, 68, 0, 0);
        nop(4);
        read(1, 71, 0, 0);
        nop(4);
        read(1, 71, 0, 0);
        nop(4);
        read(1, 71, 0, 0);
        nop(4);
        read(1, 71, 0, 0);
        nop(4);
        read(2, 52, 0, 0);
        nop(4);
        read(5, 68, 0, 0);
        nop(4);
        read(5, 68, 0, 0);
        nop(4);
        read(5, 68, 0, 0);
        nop(4);
        read(1, 71, 0, 0);
        nop(4);
        read(1, 68, 0, 0);
        nop(4);
        read(1, 68, 0, 0);
        nop(4);
        read(1, 68, 0, 0);
        nop(4);
        read(2, 52, 0, 0);
        nop(4);
        read(1, 68, 0, 0);
        nop(4);
        read(1, 68, 0, 0);
        nop(4);
        read(1, 68, 0, 0);
        nop(4);
        read(1, 68, 0, 0);
        nop(4);
        read(1, 68, 0, 0);
        nop(4);
        read(1, 69, 0, 0);
        nop(4);
        read(1, 69, 0, 0);
        nop(4);
        read(2, 52, 0, 0);
        nop(4);
        read(1, 69, 0, 0);
        nop(4);
        read(1, 69, 0, 0);
        nop(4);
        read(1, 69, 0, 0);
        nop(4);
        read(1, 69, 0, 0);
        nop(4);
        read(1, 69, 0, 0);
        nop(4);
        read(1, 69, 0, 0);
        nop(2);
        precharge(4, 0);
        nop(2);
        read(2, 52, 0, 0);
        nop(4);
        read(1, 70, 0, 0);
        nop(4);
        read(1, 70, 0, 0);
        nop(2);
        activate(4, 1883);
        nop(2);
        read(1, 70, 0, 0);
        nop(4);
        read(1, 70, 0, 0);
        nop(4);
        read(2, 57, 0, 0);
        nop(4);
        read(2, 57, 0, 0);
        nop(4);
        read(2, 57, 0, 0);
        nop(4);
        read(4, 23, 0, 0);
        nop(4);
        read(4, 23, 0, 0);
        nop(4);
        read(2, 57, 0, 0);
        nop(4);
        read(2, 57, 0, 0);
        nop(4);
        read(2, 57, 0, 0);
        nop(4);
        read(2, 57, 0, 0);
        nop(4);
        read(2, 57, 0, 0);
        nop(4);
        read(2, 63, 0, 0);
        nop(4);
        read(4, 23, 0, 0);
        nop(4);
        read(4, 23, 0, 0);
        nop(4);
        read(2, 63, 0, 0);
        nop(2);
        precharge(4, 0);
        nop(2);
        read(2, 63, 0, 0);
        nop(4);
        read(2, 63, 0, 0);
        nop(6);
        activate(4, 1883);
        nop(3);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(7, 2, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(7, 2, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(7, 2, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(11);
        precharge(3, 0);
        nop(6);
        read(4, 12, 0, 0);
        nop(2);
        precharge(1, 0);
        nop(2);
        read(4, 12, 0, 0);
        nop(2);
        activate(3, 369);
        nop(2);
        read(4, 12, 0, 0);
        nop(4);
        read(4, 12, 0, 0);
        nop(2);
        precharge(6, 0);
        nop(1);
        activate(1, 379);
        nop(1);
        read(4, 12, 0, 0);
        nop(4);
        read(3, 30, 0, 0);
        nop(2);
        precharge(4, 0);
        nop(2);
        read(3, 30, 0, 0);
        nop(2);
        activate(6, 421);
        nop(2);
        read(1, 99, 0, 0);
        nop(4);
        read(1, 99, 0, 0);
        nop(2);
        activate(4, 363);
        nop(2);
        read(1, 99, 0, 0);
        nop(4);
        read(1, 99, 0, 0);
        nop(4);
        read(3, 30, 0, 0);
        nop(4);
        read(3, 30, 0, 0);
        nop(4);
        read(3, 30, 0, 0);
        nop(4);
        read(6, 64, 0, 0);
        nop(2);
        precharge(3, 0);
        nop(2);
        read(6, 64, 0, 0);
        nop(4);
        read(1, 108, 0, 0);
        nop(4);
        read(1, 108, 0, 0);
        nop(2);
        activate(3, 2026);
        nop(2);
        read(6, 64, 0, 0);
        nop(4);
        read(6, 64, 0, 0);
        nop(4);
        read(6, 65, 0, 0);
        nop(4);
        read(6, 65, 0, 0);
        nop(4);
        read(6, 65, 0, 0);
        nop(4);
        read(1, 108, 0, 0);
        nop(4);
        read(3, 108, 0, 0);
        nop(2);
        precharge(1, 0);
        nop(2);
        read(6, 65, 0, 0);
        nop(4);
        read(6, 65, 0, 0);
        nop(4);
        read(6, 65, 0, 0);
        nop(2);
        activate(1, 1418);
        nop(2);
        read(6, 65, 0, 0);
        nop(4);
        read(6, 65, 0, 0);
        nop(9);
        write(1, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(1, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(2);
        precharge(5, 0);
        nop(2);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(4, 12, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(1, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(2);
        activate(5, 1581);
        nop(2);
        write(1, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(1, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(4, 12, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(4, 12, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(4, 12, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(11);
        precharge(1, 0);
        nop(6);
        read(5, 122, 0, 0);
        nop(4);
        read(3, 108, 0, 0);
        nop(2);
        activate(1, 379);
        nop(1);
        precharge(4, 0);
        nop(1);
        read(5, 122, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(2);
        read(5, 122, 0, 0);
        nop(4);
        read(5, 122, 0, 0);
        nop(3);
        activate(4, 1883);
        nop(1);
        read(1, 108, 0, 0);
        nop(2);
        precharge(0, 0);
        nop(2);
        read(5, 122, 0, 0);
        nop(1);
        activate(2, 377);
        nop(5);
        read(4, 12, 0, 0);
        nop(1);
        precharge(5, 0);
        nop(3);
        read(4, 12, 0, 0);
        nop(1);
        activate(0, 522);
        nop(1);
        precharge(1, 0);
        nop(2);
        read(2, 73, 0, 0);
        nop(4);
        read(2, 73, 0, 0);
        nop(1);
        activate(5, 389);
        nop(3);
        read(2, 73, 0, 0);
        nop(4);
        read(4, 12, 0, 0);
        nop(1);
        activate(1, 1418);
        nop(3);
        read(0, 62, 0, 0);
        nop(2);
        precharge(4, 0);
        nop(2);
        read(0, 62, 0, 0);
        nop(4);
        read(0, 62, 0, 0);
        nop(4);
        read(2, 73, 0, 0);
        nop(2);
        activate(4, 398);
        nop(2);
        read(0, 62, 0, 0);
        nop(9);
        read(4, 83, 0, 0);
        nop(2);
        precharge(0, 0);
        nop(2);
        read(4, 83, 0, 0);
        nop(4);
        read(4, 83, 0, 0);
        nop(4);
        read(4, 83, 0, 0);
        nop(2);
        activate(0, 1886);
        nop(7);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(5, 122, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(5, 122, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(5, 122, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(1, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(2);
        precharge(6, 0);
        nop(2);
        write(1, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(1, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(5, 122, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(2);
        activate(6, 340);
        nop(15);
        read(6, 20, 0, 0);
        nop(4);
        read(6, 20, 0, 0);
        nop(2);
        precharge(5, 0);
        nop(2);
        read(0, 9, 0, 0);
        nop(4);
        read(0, 9, 0, 0);
        nop(4);
        read(3, 108, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(1);
        activate(5, 1581);
        nop(1);
        read(6, 20, 0, 0);
        nop(2);
        precharge(3, 0);
        nop(2);
        read(6, 20, 0, 0);
        nop(4);
        read(0, 9, 0, 0);
        nop(2);
        activate(2, 503);
        nop(2);
        read(5, 122, 0, 0);
        nop(4);
        activate(3, 369);
        nop(1);
        read(5, 122, 0, 0);
        nop(4);
        read(5, 122, 0, 0);
        nop(4);
        read(0, 9, 0, 0);
        nop(4);
        read(3, 30, 0, 0);
        nop(2);
        precharge(0, 0);
        nop(2);
        read(3, 30, 0, 0);
        nop(2);
        precharge(6, 0);
        nop(2);
        read(3, 30, 0, 0);
        nop(6);
        activate(0, 384);
        nop(1);
        precharge(3, 0);
        nop(2);
        write(2, 103, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(3);
        activate(6, 340);
        nop(1);
        write(2, 103, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(0, 9, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(2);
        activate(3, 267);
        nop(2);
        write(2, 103, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(0, 9, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(0, 9, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(2);
        precharge(1, 0);
        nop(2);
        write(0, 9, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(4);
        write(2, 103, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(6);
        activate(1, 359);
        nop(11);
        read(1, 123, 0, 0);
        nop(4);
        read(3, 24, 0, 0);
        nop(4);
        read(3, 24, 0, 0);
        nop(4);
        read(6, 15, 0, 0);
        nop(4);
        read(6, 15, 0, 0);
        nop(4);
        read(6, 15, 0, 0);
        nop(4);
        read(1, 123, 0, 0);
        nop(2);
        precharge(5, 0);
        nop(2);
        read(1, 123, 0, 0);
        nop(4);
        read(3, 24, 0, 0);
        nop(4);
        read(3, 24, 0, 0);
        nop(2);
        activate(5, 409);
        nop(2);
        read(6, 15, 0, 0);
        nop(2);
        precharge(3, 0);
        nop(2);
        read(1, 123, 0, 0);
        nop(4);
        read(1, 123, 0, 0);
        nop(4);
        read(1, 123, 0, 0);
        nop(2);
        activate(3, 2026);
        nop(2);
        read(5, 73, 0, 0);
        nop(4);
        read(5, 73, 0, 0);
        nop(4);
        read(5, 73, 0, 0);
        nop(4);
        read(1, 123, 0, 0);
        nop(4);
        read(1, 123, 0, 0);
        nop(4);
        read(5, 73, 0, 0);
        nop(4);
        read(5, 77, 0, 0);
        nop(4);
        read(5, 77, 0, 0);
        nop(4);
        read(5, 77, 0, 0);
        nop(4);
        read(5, 77, 0, 0);
        nop(9);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(17);
        read(3, 108, 0, 0);
        nop(4);
        read(5, 77, 0, 0);
        nop(4);
        read(5, 77, 0, 0);
        nop(4);
        read(5, 77, 0, 0);
        nop(4);
        read(5, 77, 0, 0);
        nop(4);
        read(5, 78, 0, 0);
        nop(4);
        read(5, 78, 0, 0);
        nop(4);
        read(5, 78, 0, 0);
        nop(4);
        read(5, 78, 0, 0);
        nop(4);
        read(5, 78, 0, 0);
        nop(4);
        read(5, 78, 0, 0);
        nop(4);
        read(1, 124, 0, 0);
        nop(4);
        read(5, 78, 0, 0);
        nop(4);
        read(5, 78, 0, 0);
        nop(4);
        read(1, 124, 0, 0);
        nop(4);
        read(1, 124, 0, 0);
        nop(4);
        read(1, 124, 0, 0);
        nop(4);
        read(1, 124, 0, 0);
        nop(4);
        read(1, 124, 0, 0);
        nop(4);
        read(1, 124, 0, 0);
        nop(4);
        read(1, 124, 0, 0);
        nop(4);
        read(1, 125, 0, 0);
        nop(4);
        read(1, 125, 0, 0);
        nop(4);
        read(1, 125, 0, 0);
        nop(4);
        read(1, 125, 0, 0);
        nop(4);
        read(1, 125, 0, 0);
        nop(4);
        read(1, 125, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(2);
        read(1, 125, 0, 0);
        nop(4);
        read(1, 125, 0, 0);
        nop(6);
        activate(2, 520);
        nop(3);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(17);
        read(2, 99, 0, 0);
        nop(4);
        read(2, 99, 0, 0);
        nop(4);
        read(2, 99, 0, 0);
        nop(4);
        read(2, 99, 0, 0);
        nop(4);
        read(3, 108, 0, 0);
        nop(9);
        write(3, 108, 0, 0, 0, {{8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}, {8'h0}});
        nop(2);
        precharge(1, 0);
        nop(12);
        activate(1, 422);
        nop(9);
        precharge(3, 0);
        nop(2);
        read(1, 42, 0, 0);
        nop(4);
        read(1, 42, 0, 0);
        nop(4);
        read(1, 42, 0, 0);
        nop(2);
        activate(3, 522);
        nop(2);
        read(1, 42, 0, 0);
        nop(6);
        precharge(1, 0);
        nop(3);
        read(3, 96, 0, 0);
        nop(4);
        read(3, 96, 0, 0);
        nop(4);
        read(3, 96, 0, 0);
        nop(1);
        activate(1, 364);
        nop(1);
        precharge(6, 0);
        nop(2);
        read(3, 96, 0, 0);
        nop(4);
        read(3, 97, 0, 0);
        nop(4);
        read(3, 97, 0, 0);
        nop(2);
        activate(6, 513);
        nop(1);
        precharge(0, 0);
        nop(1);
        read(3, 97, 0, 0);
        nop(4);
        read(3, 97, 0, 0);
        nop(4);
        read(3, 103, 0, 0);
        nop(3);
        activate(0, 440);
        nop(1);
        read(3, 103, 0, 0);
        nop(4);
        read(6, 99, 0, 0);
        nop(4);
        read(6, 99, 0, 0);
        nop(4);
        read(6, 99, 0, 0);
        nop(2);
        precharge(4, 0);
        nop(2);
        read(0, 21, 0, 0);
        nop(4);
        read(3, 103, 0, 0);
        nop(4);
        read(3, 103, 0, 0);
        nop(2);
        activate(4, 407);
        nop(2);
        read(6, 99, 0, 0);
        nop(4);
        read(0, 21, 0, 0);
        nop(4);
        read(0, 21, 0, 0);
        nop(4);
        read(0, 21, 0, 0);
        nop(4);
        read(0, 21, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(2);
        read(3, 97, 0, 0);
        nop(4);
        read(3, 97, 0, 0);
        nop(4);
        read(4, 19, 0, 0);
        nop(2);
        activate(2, 407);
        nop(2);
        read(0, 21, 0, 0);
        nop(4);
        read(0, 21, 0, 0);
        nop(4);
        read(0, 21, 0, 0);
        nop(4);
        read(2, 80, 0, 0);
        nop(4);
        read(2, 80, 0, 0);
        nop(4);
        read(3, 97, 0, 0);
        nop(4);
        read(4, 19, 0, 0);
        nop(4);
        read(2, 80, 0, 0);
        nop(4);
        read(2, 80, 0, 0);
        nop(4);
        read(2, 80, 0, 0);
        nop(4);
        read(3, 97, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(2);
        read(3, 103, 0, 0);
        nop(4);
        read(3, 103, 0, 0);
        nop(2);
        precharge(6, 0);
        nop(2);
        read(3, 103, 0, 0);
        nop(2);
        activate(2, 265);
        nop(2);
        read(3, 103, 0, 0);
        nop(4);
        read(3, 98, 0, 0);
        nop(2);
        activate(6, 519);
        nop(2);
        read(3, 98, 0, 0);
        nop(4);
        read(3, 98, 0, 0);
        nop(4);
        read(4, 19, 0, 0);
        nop(4);
        read(6, 23, 0, 0);
        nop(4);
        read(6, 23, 0, 0);
        nop(4);
        read(2, 87, 0, 0);
        nop(4);
        read(2, 87, 0, 0);
        nop(4);
        read(2, 87, 0, 0);
        nop(4);
        read(2, 87, 0, 0);
        nop(4);
        read(3, 98, 0, 0);
        nop(4);
        read(4, 19, 0, 0);
        nop(4);
        read(6, 23, 0, 0);
        nop(4);
        read(6, 23, 0, 0);
        nop(4);
        read(2, 87, 0, 0);
        nop(4);
        read(3, 98, 0, 0);
        nop(2);
        precharge(2, 0);
        nop(2);
        read(3, 98, 0, 0);
        nop(4);
        read(3, 98, 0, 0);
        nop(4);
        read(4, 19, 0, 0);
        nop(2);
        activate(2, 407);
        nop(2);
        read(6, 23, 0, 0);
        nop(4);
        read(3, 98, 0, 0);
        nop(4);
        read(3, 102, 0, 0);
        nop(4);
        read(2, 80, 0, 0);
        nop(4);
        read(2, 80, 0, 0);
        nop(4);
        read(3, 102, 0, 0);
        nop(4);
        read(4, 19, 0, 0);
        nop(4);
        read(6, 23, 0, 0);
        nop(4);
        read(6, 23, 0, 0);
        nop(4);
        read(2, 80, 0, 0);
        nop(4);
        read(2, 81, 0, 0);
        nop(4);
        read(2, 81, 0, 0);
        nop(4);
        read(3, 102, 0, 0);
